** Generated for: hspiceD
** Generated on: Sep 22 16:25:40 2014
** Design library name: dummy_4_bit
** Design cell name: test_XORX2
** Design view name: schematic
.GLOBAL _gnet0 vdd! vss!
.PARAM vdd=1 v_low=0 buff_vdd=vdd v_hig=vdd


.TRAN 100e-12 10e-9 START=0.0

.OP

.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.INCLUDE "/ad/eng/users/b/o/bobzhou/Desktop/571/hw3/tech_files/45nm_HP.pm"

** Library name: NangateOpenCellLibrary
** Cell name: XOR2_X2
** View name: schematic
.subckt XOR2_X2 a b z
m_i_19 net_001 a z vss! NMOS_VTL L=50e-9 W=415e-9
m_i_24 vss! b net_001 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_19_23 net_001b a z vss! NMOS_VTL L=50e-9 W=415e-9
m_i_24_4 vss! b net_001b vss! NMOS_VTL L=50e-9 W=415e-9
m_i_0 net_000 a vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_7 vss! b net_000 vss! NMOS_VTL L=50e-9 W=415e-9
m_i_13 z net_000 vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_13_35 z net_000 vss! vss! NMOS_VTL L=50e-9 W=415e-9
m_i_30 net_002 a net_000 vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_35 vdd! b net_002 vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_41 net_003 net_000 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_41_29 net_003 net_000 vdd! vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_47 z a net_003 vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_53 net_003 b z vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_53_18 net_003 b z vdd! PMOS_VTL L=50e-9 W=630e-9
m_i_47_27 z a net_003 vdd! PMOS_VTL L=50e-9 W=630e-9
.ends XOR2_X2
** End of subcircuit definition.

** Library name: equalized_logic
** Cell name: buffer4test
** View name: schematic
.subckt buffer4test buff_vdd buff_vss input output inh_bulk_n inh_bulk_p
m1 output net14 buff_vdd inh_bulk_p pmos_vtl L=50e-9 W=1.26e-6
m3 net14 input buff_vdd inh_bulk_p pmos_vtl L=50e-9 W=1.26e-6
m0 output net14 buff_vss inh_bulk_n nmos_vtl L=50e-9 W=830e-9
m9 net14 input buff_vss inh_bulk_n nmos_vtl L=50e-9 W=830e-9
.ends buffer4test
** End of subcircuit definition.

** Library name: dummy_4_bit
** Cell name: test_XORX2
** View name: schematic
xi30 a_in b_in output XOR2_X2
f0 vpower 0 CCCS v3  1 M=1
v10 buff_vss 0 DC=0
v8 buff_vdd 0 DC=buff_vdd
v6 vss! 0 DC=0
v3 vdd! 0 DC=vdd
xi16 buff_vdd buff_vss a a_in 0 _gnet0 buffer4test
xi17 buff_vdd buff_vss b1 b_in 0 _gnet0 buffer4test
c10 vpower 0 1e-12 IC=0
c0 output 0 663e-18
v1 a 0 PWL
+ 0.000001n V_low
+ 0.100000n V_low
+ 0.100001n V_low
+ 0.200000n V_low
+ 0.200001n V_low
+ 0.300000n V_low
+ 0.300001n V_low
+ 0.400000n V_low
+ 0.400001n V_low
+ 0.500000n V_low
+ 0.500001n V_low
+ 0.600000n V_low
+ 0.600001n V_low
+ 0.700000n V_low
+ 0.700001n V_low
+ 0.800000n V_low
+ 0.800001n V_low
+ 0.900000n V_low
+ 0.900001n V_low
+ 1.000000n V_low
+ 1.000001n V_hig
+ 1.100000n V_hig
+ 1.100001n V_hig
+ 1.200000n V_hig
+ 1.200001n V_hig
+ 1.300000n V_hig
+ 1.300001n V_hig
+ 1.400000n V_hig
+ 1.400001n V_hig
+ 1.500000n V_hig
+ 1.500001n V_hig
+ 1.600000n V_hig
+ 1.600001n V_hig
+ 1.700000n V_hig
+ 1.700001n V_hig
+ 1.800000n V_hig
+ 1.800001n V_hig
+ 1.900000n V_hig
+ 1.900001n V_hig
+ 2.000000n V_hig
+ 2.000001n V_low
+ 2.100000n V_low
+ 2.100001n V_low
+ 2.200000n V_low
+ 2.200001n V_low
+ 2.300000n V_low
+ 2.300001n V_low
+ 2.400000n V_low
+ 2.400001n V_low
+ 2.500000n V_low
+ 2.500001n V_low
+ 2.600000n V_low
+ 2.600001n V_low
+ 2.700000n V_low
+ 2.700001n V_low
+ 2.800000n V_low
+ 2.800001n V_low
+ 2.900000n V_low
+ 2.900001n V_low
+ 3.000000n V_low
+ 3.000001n V_hig
+ 3.100000n V_hig
+ 3.100001n V_hig
+ 3.200000n V_hig
+ 3.200001n V_hig
+ 3.300000n V_hig
+ 3.300001n V_hig
+ 3.400000n V_hig
+ 3.400001n V_hig
+ 3.500000n V_hig
+ 3.500001n V_hig
+ 3.600000n V_hig
+ 3.600001n V_hig
+ 3.700000n V_hig
+ 3.700001n V_hig
+ 3.800000n V_hig
+ 3.800001n V_hig
+ 3.900000n V_hig
+ 3.900001n V_hig
+ 4.000000n V_hig
+ 4.000001n V_low
+ 4.100000n V_low
+ 4.100001n V_low
+ 4.200000n V_low
+ 4.200001n V_low
+ 4.300000n V_low
+ 4.300001n V_low
+ 4.400000n V_low
+ 4.400001n V_low
+ 4.500000n V_low
+ 4.500001n V_low
+ 4.600000n V_low
+ 4.600001n V_low
+ 4.700000n V_low
+ 4.700001n V_low
+ 4.800000n V_low
+ 4.800001n V_low
+ 4.900000n V_low
+ 4.900001n V_low
+ 5.000000n V_low
+ 5.000001n V_hig
+ 5.100000n V_hig
+ 5.100001n V_hig
+ 5.200000n V_hig
+ 5.200001n V_hig
+ 5.300000n V_hig
+ 5.300001n V_hig
+ 5.400000n V_hig
+ 5.400001n V_hig
+ 5.500000n V_hig
+ 5.500001n V_hig
+ 5.600000n V_hig
+ 5.600001n V_hig
+ 5.700000n V_hig
+ 5.700001n V_hig
+ 5.800000n V_hig
+ 5.800001n V_hig
+ 5.900000n V_hig
+ 5.900001n V_hig
+ 6.000000n V_hig
+ 6.000001n V_low
+ 6.100000n V_low
+ 6.100001n V_low
+ 6.200000n V_low
+ 6.200001n V_low
+ 6.300000n V_low
+ 6.300001n V_low
+ 6.400000n V_low
+ 6.400001n V_low
+ 6.500000n V_low
+ 6.500001n V_low
+ 6.600000n V_low
+ 6.600001n V_low
+ 6.700000n V_low
+ 6.700001n V_low
+ 6.800000n V_low
+ 6.800001n V_low
+ 6.900000n V_low
+ 6.900001n V_low
+ 7.000000n V_low
+ 7.000001n V_hig
+ 7.100000n V_hig
+ 7.100001n V_hig
+ 7.200000n V_hig
+ 7.200001n V_hig
+ 7.300000n V_hig
+ 7.300001n V_hig
+ 7.400000n V_hig
+ 7.400001n V_hig
+ 7.500000n V_hig
+ 7.500001n V_hig
+ 7.600000n V_hig
+ 7.600001n V_hig
+ 7.700000n V_hig
+ 7.700001n V_hig
+ 7.800000n V_hig
+ 7.800001n V_hig
+ 7.900000n V_hig
+ 7.900001n V_hig
+ 8.000000n V_hig
+ 8.000001n V_low
+ 8.100000n V_low
+ 8.100001n V_low
+ 8.200000n V_low
+ 8.200001n V_low
+ 8.300000n V_low
+ 8.300001n V_low
+ 8.400000n V_low
+ 8.400001n V_low
+ 8.500000n V_low
+ 8.500001n V_low
+ 8.600000n V_low
+ 8.600001n V_low
+ 8.700000n V_low
+ 8.700001n V_low
+ 8.800000n V_low
+ 8.800001n V_low
+ 8.900000n V_low
+ 8.900001n V_low
+ 9.000000n V_low
+ 9.000001n V_low
+ 9.100000n V_low
+ 9.100001n V_low
+ 9.200000n V_low
+ 9.200001n V_low
+ 9.300000n V_low
+ 9.300001n V_low
+ 9.400000n V_low
+ 9.400001n V_low
+ 9.500000n V_low
+ 9.500001n V_low
+ 9.600000n V_low
+ 9.600001n V_low
+ 9.700000n V_low
+ 9.700001n V_low
+ 9.800000n V_low
+ 9.800001n V_low
+ 9.900000n V_low
+ 9.900001n V_low
+ 10.000000n V_low
+ 10.000001n V_low
+ 10.100000n V_low
+ 10.100001n V_low
+ 10.200000n V_low
+ 10.200001n V_low
+ 10.300000n V_low
+ 10.300001n V_low
+ 10.400000n V_low
+ 10.400001n V_low
+ 10.500000n V_low
+ 10.500001n V_low
+ 10.600000n V_low
+ 10.600001n V_low
+ 10.700000n V_low
+ 10.700001n V_low
+ 10.800000n V_low
+ 10.800001n V_low
+ 10.900000n V_low
+ 10.900001n V_low
+ 11.000000n V_low
+ 11.000001n V_low
+ 11.100000n V_low
+ 11.100001n V_low
+ 11.200000n V_low
+ 11.200001n V_low
+ 11.300000n V_low
+ 11.300001n V_low
+ 11.400000n V_low
+ 11.400001n V_low
+ 11.500000n V_low
+ 11.500001n V_low
+ 11.600000n V_low
+ 11.600001n V_low
+ 11.700000n V_low
+ 11.700001n V_low
+ 11.800000n V_low
+ 11.800001n V_low
+ 11.900000n V_low
+ 11.900001n V_low
+ 12.000000n V_low
+ 12.000001n V_hig
+ 12.100000n V_hig
+ 12.100001n V_hig
+ 12.200000n V_hig
+ 12.200001n V_hig
+ 12.300000n V_hig
+ 12.300001n V_hig
+ 12.400000n V_hig
+ 12.400001n V_hig
+ 12.500000n V_hig
+ 12.500001n V_hig
+ 12.600000n V_hig
+ 12.600001n V_hig
+ 12.700000n V_hig
+ 12.700001n V_hig
+ 12.800000n V_hig
+ 12.800001n V_hig
+ 12.900000n V_hig
+ 12.900001n V_hig
+ 13.000000n V_hig
+ 13.000001n V_hig
+ 13.100000n V_hig
+ 13.100001n V_hig
+ 13.200000n V_hig
+ 13.200001n V_hig
+ 13.300000n V_hig
+ 13.300001n V_hig
+ 13.400000n V_hig
+ 13.400001n V_hig
+ 13.500000n V_hig
+ 13.500001n V_hig
+ 13.600000n V_hig
+ 13.600001n V_hig
+ 13.700000n V_hig
+ 13.700001n V_hig
+ 13.800000n V_hig
+ 13.800001n V_hig
+ 13.900000n V_hig
+ 13.900001n V_hig
+ 14.000000n V_hig
+ 14.000001n V_hig
+ 14.100000n V_hig
+ 14.100001n V_hig
+ 14.200000n V_hig
+ 14.200001n V_hig
+ 14.300000n V_hig
+ 14.300001n V_hig
+ 14.400000n V_hig
+ 14.400001n V_hig
+ 14.500000n V_hig
+ 14.500001n V_hig
+ 14.600000n V_hig
+ 14.600001n V_hig
+ 14.700000n V_hig
+ 14.700001n V_hig
+ 14.800000n V_hig
+ 14.800001n V_hig
+ 14.900000n V_hig
+ 14.900001n V_hig
+ 15.000000n V_hig
+ 15.000001n V_hig
+ 15.100000n V_hig
+ 15.100001n V_hig
+ 15.200000n V_hig
+ 15.200001n V_hig
+ 15.300000n V_hig
+ 15.300001n V_hig
+ 15.400000n V_hig
+ 15.400001n V_hig
+ 15.500000n V_hig
+ 15.500001n V_hig
+ 15.600000n V_hig
+ 15.600001n V_hig
+ 15.700000n V_hig
+ 15.700001n V_hig
+ 15.800000n V_hig
+ 15.800001n V_hig
+ 15.900000n V_hig
+ 15.900001n V_hig
+ 16.000000n V_hig
+ 16.000001n V_hig
+ 16.100000n V_hig
+ 16.100001n V_hig
+ 16.200000n V_hig
+ 16.200001n V_hig
+ 16.300000n V_hig
+ 16.300001n V_hig
+ 16.400000n V_hig
+ 16.400001n V_hig
+ 16.500000n V_hig
+ 16.500001n V_hig
+ 16.600000n V_hig
+ 16.600001n V_hig
+ 16.700000n V_hig
+ 16.700001n V_hig
+ 16.800000n V_hig
+ 16.800001n V_hig
+ 16.900000n V_hig
+ 16.900001n V_hig
+ 17.000000n V_hig
+ 17.000001n V_hig
+ 17.100000n V_hig
+ 17.100001n V_hig
+ 17.200000n V_hig
+ 17.200001n V_hig
+ 17.300000n V_hig
+ 17.300001n V_hig
+ 17.400000n V_hig
+ 17.400001n V_hig
+ 17.500000n V_hig
+ 17.500001n V_hig
+ 17.600000n V_hig
+ 17.600001n V_hig
+ 17.700000n V_hig
+ 17.700001n V_hig
+ 17.800000n V_hig
+ 17.800001n V_hig
+ 17.900000n V_hig
+ 17.900001n V_hig
+ 18.000000n V_hig
+ 18.000001n V_low
+ 18.100000n V_low
+ 18.100001n V_low
+ 18.200000n V_low
+ 18.200001n V_low
+ 18.300000n V_low
+ 18.300001n V_low
+ 18.400000n V_low
+ 18.400001n V_low
+ 18.500000n V_low
+ 18.500001n V_low
+ 18.600000n V_low
+ 18.600001n V_low
+ 18.700000n V_low
+ 18.700001n V_low
+ 18.800000n V_low
+ 18.800001n V_low
+ 18.900000n V_low
+ 18.900001n V_low
+ 19.000000n V_low
+ 19.000001n V_low
+ 19.100000n V_low
+ 19.100001n V_low
+ 19.200000n V_low
+ 19.200001n V_low
+ 19.300000n V_low
+ 19.300001n V_low
+ 19.400000n V_low
+ 19.400001n V_low
+ 19.500000n V_low
+ 19.500001n V_low
+ 19.600000n V_low
+ 19.600001n V_low
+ 19.700000n V_low
+ 19.700001n V_low
+ 19.800000n V_low
+ 19.800001n V_low
+ 19.900000n V_low
+ 19.900001n V_low
+ 20.000000n V_low
+ 20.000001n V_low
+ 20.100000n V_low
+ 20.100001n V_low
+ 20.200000n V_low
+ 20.200001n V_low
+ 20.300000n V_low
+ 20.300001n V_low
+ 20.400000n V_low
+ 20.400001n V_low
+ 20.500000n V_low
+ 20.500001n V_low
+ 20.600000n V_low
+ 20.600001n V_low
+ 20.700000n V_low
+ 20.700001n V_low
+ 20.800000n V_low
+ 20.800001n V_low
+ 20.900000n V_low
+ 20.900001n V_low
+ 21.000000n V_low
+ 21.000001n V_hig
+ 21.100000n V_hig
+ 21.100001n V_hig
+ 21.200000n V_hig
+ 21.200001n V_hig
+ 21.300000n V_hig
+ 21.300001n V_hig
+ 21.400000n V_hig
+ 21.400001n V_hig
+ 21.500000n V_hig
+ 21.500001n V_hig
+ 21.600000n V_hig
+ 21.600001n V_hig
+ 21.700000n V_hig
+ 21.700001n V_hig
+ 21.800000n V_hig
+ 21.800001n V_hig
+ 21.900000n V_hig
+ 21.900001n V_hig
+ 22.000000n V_hig
+ 22.000001n V_low
+ 22.100000n V_low
+ 22.100001n V_low
+ 22.200000n V_low
+ 22.200001n V_low
+ 22.300000n V_low
+ 22.300001n V_low
+ 22.400000n V_low
+ 22.400001n V_low
+ 22.500000n V_low
+ 22.500001n V_low
+ 22.600000n V_low
+ 22.600001n V_low
+ 22.700000n V_low
+ 22.700001n V_low
+ 22.800000n V_low
+ 22.800001n V_low
+ 22.900000n V_low
+ 22.900001n V_low
+ 23.000000n V_low
+ 23.000001n V_hig
+ 23.100000n V_hig
+ 23.100001n V_hig
+ 23.200000n V_hig
+ 23.200001n V_hig
+ 23.300000n V_hig
+ 23.300001n V_hig
+ 23.400000n V_hig
+ 23.400001n V_hig
+ 23.500000n V_hig
+ 23.500001n V_hig
+ 23.600000n V_hig
+ 23.600001n V_hig
+ 23.700000n V_hig
+ 23.700001n V_hig
+ 23.800000n V_hig
+ 23.800001n V_hig
+ 23.900000n V_hig
+ 23.900001n V_hig
+ 24.000000n V_hig
+ 24.000001n V_hig
+ 24.100000n V_hig
+ 24.100001n V_hig
+ 24.200000n V_hig
+ 24.200001n V_hig
+ 24.300000n V_hig
+ 24.300001n V_hig
+ 24.400000n V_hig
+ 24.400001n V_hig
+ 24.500000n V_hig
+ 24.500001n V_hig
+ 24.600000n V_hig
+ 24.600001n V_hig
+ 24.700000n V_hig
+ 24.700001n V_hig
+ 24.800000n V_hig
+ 24.800001n V_hig
+ 24.900000n V_hig
+ 24.900001n V_hig
+ 25.000000n V_hig
+ 25.000001n V_hig
+ 25.100000n V_hig
+ 25.100001n V_hig
+ 25.200000n V_hig
+ 25.200001n V_hig
+ 25.300000n V_hig
+ 25.300001n V_hig
+ 25.400000n V_hig
+ 25.400001n V_hig
+ 25.500000n V_hig
+ 25.500001n V_hig
+ 25.600000n V_hig
+ 25.600001n V_hig
+ 25.700000n V_hig
+ 25.700001n V_hig
+ 25.800000n V_hig
+ 25.800001n V_hig
+ 25.900000n V_hig
+ 25.900001n V_hig
+ 26.000000n V_hig
+ 26.000001n V_hig
+ 26.100000n V_hig
+ 26.100001n V_hig
+ 26.200000n V_hig
+ 26.200001n V_hig
+ 26.300000n V_hig
+ 26.300001n V_hig
+ 26.400000n V_hig
+ 26.400001n V_hig
+ 26.500000n V_hig
+ 26.500001n V_hig
+ 26.600000n V_hig
+ 26.600001n V_hig
+ 26.700000n V_hig
+ 26.700001n V_hig
+ 26.800000n V_hig
+ 26.800001n V_hig
+ 26.900000n V_hig
+ 26.900001n V_hig
+ 27.000000n V_hig
+ 27.000001n V_low
+ 27.100000n V_low
+ 27.100001n V_low
+ 27.200000n V_low
+ 27.200001n V_low
+ 27.300000n V_low
+ 27.300001n V_low
+ 27.400000n V_low
+ 27.400001n V_low
+ 27.500000n V_low
+ 27.500001n V_low
+ 27.600000n V_low
+ 27.600001n V_low
+ 27.700000n V_low
+ 27.700001n V_low
+ 27.800000n V_low
+ 27.800001n V_low
+ 27.900000n V_low
+ 27.900001n V_low
+ 28.000000n V_low
+ 28.000001n V_low
+ 28.100000n V_low
+ 28.100001n V_low
+ 28.200000n V_low
+ 28.200001n V_low
+ 28.300000n V_low
+ 28.300001n V_low
+ 28.400000n V_low
+ 28.400001n V_low
+ 28.500000n V_low
+ 28.500001n V_low
+ 28.600000n V_low
+ 28.600001n V_low
+ 28.700000n V_low
+ 28.700001n V_low
+ 28.800000n V_low
+ 28.800001n V_low
+ 28.900000n V_low
+ 28.900001n V_low
+ 29.000000n V_low
+ 29.000001n V_hig
+ 29.100000n V_hig
+ 29.100001n V_hig
+ 29.200000n V_hig
+ 29.200001n V_hig
+ 29.300000n V_hig
+ 29.300001n V_hig
+ 29.400000n V_hig
+ 29.400001n V_hig
+ 29.500000n V_hig
+ 29.500001n V_hig
+ 29.600000n V_hig
+ 29.600001n V_hig
+ 29.700000n V_hig
+ 29.700001n V_hig
+ 29.800000n V_hig
+ 29.800001n V_hig
+ 29.900000n V_hig
+ 29.900001n V_hig
+ 30.000000n V_hig
+ 30.000001n V_hig
+ 30.100000n V_hig
+ 30.100001n V_hig
+ 30.200000n V_hig
+ 30.200001n V_hig
+ 30.300000n V_hig
+ 30.300001n V_hig
+ 30.400000n V_hig
+ 30.400001n V_hig
+ 30.500000n V_hig
+ 30.500001n V_hig
+ 30.600000n V_hig
+ 30.600001n V_hig
+ 30.700000n V_hig
+ 30.700001n V_hig
+ 30.800000n V_hig
+ 30.800001n V_hig
+ 30.900000n V_hig
+ 30.900001n V_hig
+ 31.000000n V_hig
+ 31.000001n V_low
+ 31.100000n V_low
+ 31.100001n V_low
+ 31.200000n V_low
+ 31.200001n V_low
+ 31.300000n V_low
+ 31.300001n V_low
+ 31.400000n V_low
+ 31.400001n V_low
+ 31.500000n V_low
+ 31.500001n V_low
+ 31.600000n V_low
+ 31.600001n V_low
+ 31.700000n V_low
+ 31.700001n V_low
+ 31.800000n V_low
+ 31.800001n V_low
+ 31.900000n V_low
+ 31.900001n V_low
+ 32.000000n V_low
+ 32.000001n V_low
+ 32.100000n V_low
+ 32.100001n V_low
+ 32.200000n V_low
+ 32.200001n V_low
+ 32.300000n V_low
+ 32.300001n V_low
+ 32.400000n V_low
+ 32.400001n V_low
+ 32.500000n V_low
+ 32.500001n V_low
+ 32.600000n V_low
+ 32.600001n V_low
+ 32.700000n V_low
+ 32.700001n V_low
+ 32.800000n V_low
+ 32.800001n V_low
+ 32.900000n V_low
+ 32.900001n V_low
+ 33.000000n V_low
+ 33.000001n V_low
+ 33.100000n V_low
+ 33.100001n V_low
+ 33.200000n V_low
+ 33.200001n V_low
+ 33.300000n V_low
+ 33.300001n V_low
+ 33.400000n V_low
+ 33.400001n V_low
+ 33.500000n V_low
+ 33.500001n V_low
+ 33.600000n V_low
+ 33.600001n V_low
+ 33.700000n V_low
+ 33.700001n V_low
+ 33.800000n V_low
+ 33.800001n V_low
+ 33.900000n V_low
+ 33.900001n V_low
+ 34.000000n V_low
+ 34.000001n V_low
+ 34.100000n V_low
+ 34.100001n V_low
+ 34.200000n V_low
+ 34.200001n V_low
+ 34.300000n V_low
+ 34.300001n V_low
+ 34.400000n V_low
+ 34.400001n V_low
+ 34.500000n V_low
+ 34.500001n V_low
+ 34.600000n V_low
+ 34.600001n V_low
+ 34.700000n V_low
+ 34.700001n V_low
+ 34.800000n V_low
+ 34.800001n V_low
+ 34.900000n V_low
+ 34.900001n V_low
+ 35.000000n V_low
+ 35.000001n V_low
+ 35.100000n V_low
+ 35.100001n V_low
+ 35.200000n V_low
+ 35.200001n V_low
+ 35.300000n V_low
+ 35.300001n V_low
+ 35.400000n V_low
+ 35.400001n V_low
+ 35.500000n V_low
+ 35.500001n V_low
+ 35.600000n V_low
+ 35.600001n V_low
+ 35.700000n V_low
+ 35.700001n V_low
+ 35.800000n V_low
+ 35.800001n V_low
+ 35.900000n V_low
+ 35.900001n V_low
+ 36.000000n V_low
+ 36.000001n V_low
+ 36.100000n V_low
+ 36.100001n V_low
+ 36.200000n V_low
+ 36.200001n V_low
+ 36.300000n V_low
+ 36.300001n V_low
+ 36.400000n V_low
+ 36.400001n V_low
+ 36.500000n V_low
+ 36.500001n V_low
+ 36.600000n V_low
+ 36.600001n V_low
+ 36.700000n V_low
+ 36.700001n V_low
+ 36.800000n V_low
+ 36.800001n V_low
+ 36.900000n V_low
+ 36.900001n V_low
+ 37.000000n V_low
+ 37.000001n V_hig
+ 37.100000n V_hig
+ 37.100001n V_hig
+ 37.200000n V_hig
+ 37.200001n V_hig
+ 37.300000n V_hig
+ 37.300001n V_hig
+ 37.400000n V_hig
+ 37.400001n V_hig
+ 37.500000n V_hig
+ 37.500001n V_hig
+ 37.600000n V_hig
+ 37.600001n V_hig
+ 37.700000n V_hig
+ 37.700001n V_hig
+ 37.800000n V_hig
+ 37.800001n V_hig
+ 37.900000n V_hig
+ 37.900001n V_hig
+ 38.000000n V_hig
+ 38.000001n V_low
+ 38.100000n V_low
+ 38.100001n V_low
+ 38.200000n V_low
+ 38.200001n V_low
+ 38.300000n V_low
+ 38.300001n V_low
+ 38.400000n V_low
+ 38.400001n V_low
+ 38.500000n V_low
+ 38.500001n V_low
+ 38.600000n V_low
+ 38.600001n V_low
+ 38.700000n V_low
+ 38.700001n V_low
+ 38.800000n V_low
+ 38.800001n V_low
+ 38.900000n V_low
+ 38.900001n V_low
+ 39.000000n V_low
+ 39.000001n V_low
+ 39.100000n V_low
+ 39.100001n V_low
+ 39.200000n V_low
+ 39.200001n V_low
+ 39.300000n V_low
+ 39.300001n V_low
+ 39.400000n V_low
+ 39.400001n V_low
+ 39.500000n V_low
+ 39.500001n V_low
+ 39.600000n V_low
+ 39.600001n V_low
+ 39.700000n V_low
+ 39.700001n V_low
+ 39.800000n V_low
+ 39.800001n V_low
+ 39.900000n V_low
+ 39.900001n V_low
+ 40.000000n V_low
+ 40.000001n V_low
+ 40.100000n V_low
+ 40.100001n V_low
+ 40.200000n V_low
+ 40.200001n V_low
+ 40.300000n V_low
+ 40.300001n V_low
+ 40.400000n V_low
+ 40.400001n V_low
+ 40.500000n V_low
+ 40.500001n V_low
+ 40.600000n V_low
+ 40.600001n V_low
+ 40.700000n V_low
+ 40.700001n V_low
+ 40.800000n V_low
+ 40.800001n V_low
+ 40.900000n V_low
+ 40.900001n V_low
+ 41.000000n V_low
+ 41.000001n V_hig
+ 41.100000n V_hig
+ 41.100001n V_hig
+ 41.200000n V_hig
+ 41.200001n V_hig
+ 41.300000n V_hig
+ 41.300001n V_hig
+ 41.400000n V_hig
+ 41.400001n V_hig
+ 41.500000n V_hig
+ 41.500001n V_hig
+ 41.600000n V_hig
+ 41.600001n V_hig
+ 41.700000n V_hig
+ 41.700001n V_hig
+ 41.800000n V_hig
+ 41.800001n V_hig
+ 41.900000n V_hig
+ 41.900001n V_hig
+ 42.000000n V_hig
+ 42.000001n V_hig
+ 42.100000n V_hig
+ 42.100001n V_hig
+ 42.200000n V_hig
+ 42.200001n V_hig
+ 42.300000n V_hig
+ 42.300001n V_hig
+ 42.400000n V_hig
+ 42.400001n V_hig
+ 42.500000n V_hig
+ 42.500001n V_hig
+ 42.600000n V_hig
+ 42.600001n V_hig
+ 42.700000n V_hig
+ 42.700001n V_hig
+ 42.800000n V_hig
+ 42.800001n V_hig
+ 42.900000n V_hig
+ 42.900001n V_hig
+ 43.000000n V_hig
+ 43.000001n V_low
+ 43.100000n V_low
+ 43.100001n V_low
+ 43.200000n V_low
+ 43.200001n V_low
+ 43.300000n V_low
+ 43.300001n V_low
+ 43.400000n V_low
+ 43.400001n V_low
+ 43.500000n V_low
+ 43.500001n V_low
+ 43.600000n V_low
+ 43.600001n V_low
+ 43.700000n V_low
+ 43.700001n V_low
+ 43.800000n V_low
+ 43.800001n V_low
+ 43.900000n V_low
+ 43.900001n V_low
+ 44.000000n V_low
+ 44.000001n V_low
+ 44.100000n V_low
+ 44.100001n V_low
+ 44.200000n V_low
+ 44.200001n V_low
+ 44.300000n V_low
+ 44.300001n V_low
+ 44.400000n V_low
+ 44.400001n V_low
+ 44.500000n V_low
+ 44.500001n V_low
+ 44.600000n V_low
+ 44.600001n V_low
+ 44.700000n V_low
+ 44.700001n V_low
+ 44.800000n V_low
+ 44.800001n V_low
+ 44.900000n V_low
+ 44.900001n V_low
+ 45.000000n V_low
+ 45.000001n V_low
+ 45.100000n V_low
+ 45.100001n V_low
+ 45.200000n V_low
+ 45.200001n V_low
+ 45.300000n V_low
+ 45.300001n V_low
+ 45.400000n V_low
+ 45.400001n V_low
+ 45.500000n V_low
+ 45.500001n V_low
+ 45.600000n V_low
+ 45.600001n V_low
+ 45.700000n V_low
+ 45.700001n V_low
+ 45.800000n V_low
+ 45.800001n V_low
+ 45.900000n V_low
+ 45.900001n V_low
+ 46.000000n V_low
+ 46.000001n V_hig
+ 46.100000n V_hig
+ 46.100001n V_hig
+ 46.200000n V_hig
+ 46.200001n V_hig
+ 46.300000n V_hig
+ 46.300001n V_hig
+ 46.400000n V_hig
+ 46.400001n V_hig
+ 46.500000n V_hig
+ 46.500001n V_hig
+ 46.600000n V_hig
+ 46.600001n V_hig
+ 46.700000n V_hig
+ 46.700001n V_hig
+ 46.800000n V_hig
+ 46.800001n V_hig
+ 46.900000n V_hig
+ 46.900001n V_hig
+ 47.000000n V_hig
+ 47.000001n V_hig
+ 47.100000n V_hig
+ 47.100001n V_hig
+ 47.200000n V_hig
+ 47.200001n V_hig
+ 47.300000n V_hig
+ 47.300001n V_hig
+ 47.400000n V_hig
+ 47.400001n V_hig
+ 47.500000n V_hig
+ 47.500001n V_hig
+ 47.600000n V_hig
+ 47.600001n V_hig
+ 47.700000n V_hig
+ 47.700001n V_hig
+ 47.800000n V_hig
+ 47.800001n V_hig
+ 47.900000n V_hig
+ 47.900001n V_hig
+ 48.000000n V_hig
+ 48.000001n V_low
+ 48.100000n V_low
+ 48.100001n V_low
+ 48.200000n V_low
+ 48.200001n V_low
+ 48.300000n V_low
+ 48.300001n V_low
+ 48.400000n V_low
+ 48.400001n V_low
+ 48.500000n V_low
+ 48.500001n V_low
+ 48.600000n V_low
+ 48.600001n V_low
+ 48.700000n V_low
+ 48.700001n V_low
+ 48.800000n V_low
+ 48.800001n V_low
+ 48.900000n V_low
+ 48.900001n V_low
+ 49.000000n V_low
+ 49.000001n V_hig
+ 49.100000n V_hig
+ 49.100001n V_hig
+ 49.200000n V_hig
+ 49.200001n V_hig
+ 49.300000n V_hig
+ 49.300001n V_hig
+ 49.400000n V_hig
+ 49.400001n V_hig
+ 49.500000n V_hig
+ 49.500001n V_hig
+ 49.600000n V_hig
+ 49.600001n V_hig
+ 49.700000n V_hig
+ 49.700001n V_hig
+ 49.800000n V_hig
+ 49.800001n V_hig
+ 49.900000n V_hig
+ 49.900001n V_hig
+ 50.000000n V_hig
+ 50.000001n V_low
+ 50.100000n V_low
+ 50.100001n V_low
+ 50.200000n V_low
+ 50.200001n V_low
+ 50.300000n V_low
+ 50.300001n V_low
+ 50.400000n V_low
+ 50.400001n V_low
+ 50.500000n V_low
+ 50.500001n V_low
+ 50.600000n V_low
+ 50.600001n V_low
+ 50.700000n V_low
+ 50.700001n V_low
+ 50.800000n V_low
+ 50.800001n V_low
+ 50.900000n V_low
+ 50.900001n V_low
+ 51.000000n V_low
+ 51.000001n V_hig
+ 51.100000n V_hig
+ 51.100001n V_hig
+ 51.200000n V_hig
+ 51.200001n V_hig
+ 51.300000n V_hig
+ 51.300001n V_hig
+ 51.400000n V_hig
+ 51.400001n V_hig
+ 51.500000n V_hig
+ 51.500001n V_hig
+ 51.600000n V_hig
+ 51.600001n V_hig
+ 51.700000n V_hig
+ 51.700001n V_hig
+ 51.800000n V_hig
+ 51.800001n V_hig
+ 51.900000n V_hig
+ 51.900001n V_hig
+ 52.000000n V_hig
+ 52.000001n V_hig
+ 52.100000n V_hig
+ 52.100001n V_hig
+ 52.200000n V_hig
+ 52.200001n V_hig
+ 52.300000n V_hig
+ 52.300001n V_hig
+ 52.400000n V_hig
+ 52.400001n V_hig
+ 52.500000n V_hig
+ 52.500001n V_hig
+ 52.600000n V_hig
+ 52.600001n V_hig
+ 52.700000n V_hig
+ 52.700001n V_hig
+ 52.800000n V_hig
+ 52.800001n V_hig
+ 52.900000n V_hig
+ 52.900001n V_hig
+ 53.000000n V_hig
+ 53.000001n V_low
+ 53.100000n V_low
+ 53.100001n V_low
+ 53.200000n V_low
+ 53.200001n V_low
+ 53.300000n V_low
+ 53.300001n V_low
+ 53.400000n V_low
+ 53.400001n V_low
+ 53.500000n V_low
+ 53.500001n V_low
+ 53.600000n V_low
+ 53.600001n V_low
+ 53.700000n V_low
+ 53.700001n V_low
+ 53.800000n V_low
+ 53.800001n V_low
+ 53.900000n V_low
+ 53.900001n V_low
+ 54.000000n V_low
+ 54.000001n V_low
+ 54.100000n V_low
+ 54.100001n V_low
+ 54.200000n V_low
+ 54.200001n V_low
+ 54.300000n V_low
+ 54.300001n V_low
+ 54.400000n V_low
+ 54.400001n V_low
+ 54.500000n V_low
+ 54.500001n V_low
+ 54.600000n V_low
+ 54.600001n V_low
+ 54.700000n V_low
+ 54.700001n V_low
+ 54.800000n V_low
+ 54.800001n V_low
+ 54.900000n V_low
+ 54.900001n V_low
+ 55.000000n V_low
+ 55.000001n V_hig
+ 55.100000n V_hig
+ 55.100001n V_hig
+ 55.200000n V_hig
+ 55.200001n V_hig
+ 55.300000n V_hig
+ 55.300001n V_hig
+ 55.400000n V_hig
+ 55.400001n V_hig
+ 55.500000n V_hig
+ 55.500001n V_hig
+ 55.600000n V_hig
+ 55.600001n V_hig
+ 55.700000n V_hig
+ 55.700001n V_hig
+ 55.800000n V_hig
+ 55.800001n V_hig
+ 55.900000n V_hig
+ 55.900001n V_hig
+ 56.000000n V_hig
+ 56.000001n V_low
+ 56.100000n V_low
+ 56.100001n V_low
+ 56.200000n V_low
+ 56.200001n V_low
+ 56.300000n V_low
+ 56.300001n V_low
+ 56.400000n V_low
+ 56.400001n V_low
+ 56.500000n V_low
+ 56.500001n V_low
+ 56.600000n V_low
+ 56.600001n V_low
+ 56.700000n V_low
+ 56.700001n V_low
+ 56.800000n V_low
+ 56.800001n V_low
+ 56.900000n V_low
+ 56.900001n V_low
+ 57.000000n V_low
+ 57.000001n V_low
+ 57.100000n V_low
+ 57.100001n V_low
+ 57.200000n V_low
+ 57.200001n V_low
+ 57.300000n V_low
+ 57.300001n V_low
+ 57.400000n V_low
+ 57.400001n V_low
+ 57.500000n V_low
+ 57.500001n V_low
+ 57.600000n V_low
+ 57.600001n V_low
+ 57.700000n V_low
+ 57.700001n V_low
+ 57.800000n V_low
+ 57.800001n V_low
+ 57.900000n V_low
+ 57.900001n V_low
+ 58.000000n V_low
+ 58.000001n V_hig
+ 58.100000n V_hig
+ 58.100001n V_hig
+ 58.200000n V_hig
+ 58.200001n V_hig
+ 58.300000n V_hig
+ 58.300001n V_hig
+ 58.400000n V_hig
+ 58.400001n V_hig
+ 58.500000n V_hig
+ 58.500001n V_hig
+ 58.600000n V_hig
+ 58.600001n V_hig
+ 58.700000n V_hig
+ 58.700001n V_hig
+ 58.800000n V_hig
+ 58.800001n V_hig
+ 58.900000n V_hig
+ 58.900001n V_hig
+ 59.000000n V_hig
+ 59.000001n V_low
+ 59.100000n V_low
+ 59.100001n V_low
+ 59.200000n V_low
+ 59.200001n V_low
+ 59.300000n V_low
+ 59.300001n V_low
+ 59.400000n V_low
+ 59.400001n V_low
+ 59.500000n V_low
+ 59.500001n V_low
+ 59.600000n V_low
+ 59.600001n V_low
+ 59.700000n V_low
+ 59.700001n V_low
+ 59.800000n V_low
+ 59.800001n V_low
+ 59.900000n V_low
+ 59.900001n V_low
+ 60.000000n V_low
+ 60.000001n V_low
+ 60.100000n V_low
+ 60.100001n V_low
+ 60.200000n V_low
+ 60.200001n V_low
+ 60.300000n V_low
+ 60.300001n V_low
+ 60.400000n V_low
+ 60.400001n V_low
+ 60.500000n V_low
+ 60.500001n V_low
+ 60.600000n V_low
+ 60.600001n V_low
+ 60.700000n V_low
+ 60.700001n V_low
+ 60.800000n V_low
+ 60.800001n V_low
+ 60.900000n V_low
+ 60.900001n V_low
+ 61.000000n V_low
+ 61.000001n V_hig
+ 61.100000n V_hig
+ 61.100001n V_hig
+ 61.200000n V_hig
+ 61.200001n V_hig
+ 61.300000n V_hig
+ 61.300001n V_hig
+ 61.400000n V_hig
+ 61.400001n V_hig
+ 61.500000n V_hig
+ 61.500001n V_hig
+ 61.600000n V_hig
+ 61.600001n V_hig
+ 61.700000n V_hig
+ 61.700001n V_hig
+ 61.800000n V_hig
+ 61.800001n V_hig
+ 61.900000n V_hig
+ 61.900001n V_hig
+ 62.000000n V_hig
+ 62.000001n V_low
+ 62.100000n V_low
+ 62.100001n V_low
+ 62.200000n V_low
+ 62.200001n V_low
+ 62.300000n V_low
+ 62.300001n V_low
+ 62.400000n V_low
+ 62.400001n V_low
+ 62.500000n V_low
+ 62.500001n V_low
+ 62.600000n V_low
+ 62.600001n V_low
+ 62.700000n V_low
+ 62.700001n V_low
+ 62.800000n V_low
+ 62.800001n V_low
+ 62.900000n V_low
+ 62.900001n V_low
+ 63.000000n V_low
+ 63.000001n V_low
+ 63.100000n V_low
+ 63.100001n V_low
+ 63.200000n V_low
+ 63.200001n V_low
+ 63.300000n V_low
+ 63.300001n V_low
+ 63.400000n V_low
+ 63.400001n V_low
+ 63.500000n V_low
+ 63.500001n V_low
+ 63.600000n V_low
+ 63.600001n V_low
+ 63.700000n V_low
+ 63.700001n V_low
+ 63.800000n V_low
+ 63.800001n V_low
+ 63.900000n V_low
+ 63.900001n V_low
+ 64.000000n V_low
+ 64.000001n V_hig
+ 64.100000n V_hig
+ 64.100001n V_hig
+ 64.200000n V_hig
+ 64.200001n V_hig
+ 64.300000n V_hig
+ 64.300001n V_hig
+ 64.400000n V_hig
+ 64.400001n V_hig
+ 64.500000n V_hig
+ 64.500001n V_hig
+ 64.600000n V_hig
+ 64.600001n V_hig
+ 64.700000n V_hig
+ 64.700001n V_hig
+ 64.800000n V_hig
+ 64.800001n V_hig
+ 64.900000n V_hig
+ 64.900001n V_hig
+ 65.000000n V_hig
+ 65.000001n V_hig
+ 65.100000n V_hig
+ 65.100001n V_hig
+ 65.200000n V_hig
+ 65.200001n V_hig
+ 65.300000n V_hig
+ 65.300001n V_hig
+ 65.400000n V_hig
+ 65.400001n V_hig
+ 65.500000n V_hig
+ 65.500001n V_hig
+ 65.600000n V_hig
+ 65.600001n V_hig
+ 65.700000n V_hig
+ 65.700001n V_hig
+ 65.800000n V_hig
+ 65.800001n V_hig
+ 65.900000n V_hig
+ 65.900001n V_hig
+ 66.000000n V_hig
+ 66.000001n V_low
+ 66.100000n V_low
+ 66.100001n V_low
+ 66.200000n V_low
+ 66.200001n V_low
+ 66.300000n V_low
+ 66.300001n V_low
+ 66.400000n V_low
+ 66.400001n V_low
+ 66.500000n V_low
+ 66.500001n V_low
+ 66.600000n V_low
+ 66.600001n V_low
+ 66.700000n V_low
+ 66.700001n V_low
+ 66.800000n V_low
+ 66.800001n V_low
+ 66.900000n V_low
+ 66.900001n V_low
+ 67.000000n V_low
+ 67.000001n V_hig
+ 67.100000n V_hig
+ 67.100001n V_hig
+ 67.200000n V_hig
+ 67.200001n V_hig
+ 67.300000n V_hig
+ 67.300001n V_hig
+ 67.400000n V_hig
+ 67.400001n V_hig
+ 67.500000n V_hig
+ 67.500001n V_hig
+ 67.600000n V_hig
+ 67.600001n V_hig
+ 67.700000n V_hig
+ 67.700001n V_hig
+ 67.800000n V_hig
+ 67.800001n V_hig
+ 67.900000n V_hig
+ 67.900001n V_hig
+ 68.000000n V_hig
+ 68.000001n V_low
+ 68.100000n V_low
+ 68.100001n V_low
+ 68.200000n V_low
+ 68.200001n V_low
+ 68.300000n V_low
+ 68.300001n V_low
+ 68.400000n V_low
+ 68.400001n V_low
+ 68.500000n V_low
+ 68.500001n V_low
+ 68.600000n V_low
+ 68.600001n V_low
+ 68.700000n V_low
+ 68.700001n V_low
+ 68.800000n V_low
+ 68.800001n V_low
+ 68.900000n V_low
+ 68.900001n V_low
+ 69.000000n V_low
+ 69.000001n V_low
+ 69.100000n V_low
+ 69.100001n V_low
+ 69.200000n V_low
+ 69.200001n V_low
+ 69.300000n V_low
+ 69.300001n V_low
+ 69.400000n V_low
+ 69.400001n V_low
+ 69.500000n V_low
+ 69.500001n V_low
+ 69.600000n V_low
+ 69.600001n V_low
+ 69.700000n V_low
+ 69.700001n V_low
+ 69.800000n V_low
+ 69.800001n V_low
+ 69.900000n V_low
+ 69.900001n V_low
+ 70.000000n V_low
+ 70.000001n V_hig
+ 70.100000n V_hig
+ 70.100001n V_hig
+ 70.200000n V_hig
+ 70.200001n V_hig
+ 70.300000n V_hig
+ 70.300001n V_hig
+ 70.400000n V_hig
+ 70.400001n V_hig
+ 70.500000n V_hig
+ 70.500001n V_hig
+ 70.600000n V_hig
+ 70.600001n V_hig
+ 70.700000n V_hig
+ 70.700001n V_hig
+ 70.800000n V_hig
+ 70.800001n V_hig
+ 70.900000n V_hig
+ 70.900001n V_hig
+ 71.000000n V_hig
+ 71.000001n V_low
+ 71.100000n V_low
+ 71.100001n V_low
+ 71.200000n V_low
+ 71.200001n V_low
+ 71.300000n V_low
+ 71.300001n V_low
+ 71.400000n V_low
+ 71.400001n V_low
+ 71.500000n V_low
+ 71.500001n V_low
+ 71.600000n V_low
+ 71.600001n V_low
+ 71.700000n V_low
+ 71.700001n V_low
+ 71.800000n V_low
+ 71.800001n V_low
+ 71.900000n V_low
+ 71.900001n V_low
+ 72.000000n V_low
+ 72.000001n V_hig
+ 72.100000n V_hig
+ 72.100001n V_hig
+ 72.200000n V_hig
+ 72.200001n V_hig
+ 72.300000n V_hig
+ 72.300001n V_hig
+ 72.400000n V_hig
+ 72.400001n V_hig
+ 72.500000n V_hig
+ 72.500001n V_hig
+ 72.600000n V_hig
+ 72.600001n V_hig
+ 72.700000n V_hig
+ 72.700001n V_hig
+ 72.800000n V_hig
+ 72.800001n V_hig
+ 72.900000n V_hig
+ 72.900001n V_hig
+ 73.000000n V_hig
+ 73.000001n V_hig
+ 73.100000n V_hig
+ 73.100001n V_hig
+ 73.200000n V_hig
+ 73.200001n V_hig
+ 73.300000n V_hig
+ 73.300001n V_hig
+ 73.400000n V_hig
+ 73.400001n V_hig
+ 73.500000n V_hig
+ 73.500001n V_hig
+ 73.600000n V_hig
+ 73.600001n V_hig
+ 73.700000n V_hig
+ 73.700001n V_hig
+ 73.800000n V_hig
+ 73.800001n V_hig
+ 73.900000n V_hig
+ 73.900001n V_hig
+ 74.000000n V_hig
+ 74.000001n V_low
+ 74.100000n V_low
+ 74.100001n V_low
+ 74.200000n V_low
+ 74.200001n V_low
+ 74.300000n V_low
+ 74.300001n V_low
+ 74.400000n V_low
+ 74.400001n V_low
+ 74.500000n V_low
+ 74.500001n V_low
+ 74.600000n V_low
+ 74.600001n V_low
+ 74.700000n V_low
+ 74.700001n V_low
+ 74.800000n V_low
+ 74.800001n V_low
+ 74.900000n V_low
+ 74.900001n V_low
+ 75.000000n V_low
+ 75.000001n V_low
+ 75.100000n V_low
+ 75.100001n V_low
+ 75.200000n V_low
+ 75.200001n V_low
+ 75.300000n V_low
+ 75.300001n V_low
+ 75.400000n V_low
+ 75.400001n V_low
+ 75.500000n V_low
+ 75.500001n V_low
+ 75.600000n V_low
+ 75.600001n V_low
+ 75.700000n V_low
+ 75.700001n V_low
+ 75.800000n V_low
+ 75.800001n V_low
+ 75.900000n V_low
+ 75.900001n V_low
+ 76.000000n V_low
+ 76.000001n V_low
+ 76.100000n V_low
+ 76.100001n V_low
+ 76.200000n V_low
+ 76.200001n V_low
+ 76.300000n V_low
+ 76.300001n V_low
+ 76.400000n V_low
+ 76.400001n V_low
+ 76.500000n V_low
+ 76.500001n V_low
+ 76.600000n V_low
+ 76.600001n V_low
+ 76.700000n V_low
+ 76.700001n V_low
+ 76.800000n V_low
+ 76.800001n V_low
+ 76.900000n V_low
+ 76.900001n V_low
+ 77.000000n V_low
+ 77.000001n V_low
+ 77.100000n V_low
+ 77.100001n V_low
+ 77.200000n V_low
+ 77.200001n V_low
+ 77.300000n V_low
+ 77.300001n V_low
+ 77.400000n V_low
+ 77.400001n V_low
+ 77.500000n V_low
+ 77.500001n V_low
+ 77.600000n V_low
+ 77.600001n V_low
+ 77.700000n V_low
+ 77.700001n V_low
+ 77.800000n V_low
+ 77.800001n V_low
+ 77.900000n V_low
+ 77.900001n V_low
+ 78.000000n V_low
+ 78.000001n V_hig
+ 78.100000n V_hig
+ 78.100001n V_hig
+ 78.200000n V_hig
+ 78.200001n V_hig
+ 78.300000n V_hig
+ 78.300001n V_hig
+ 78.400000n V_hig
+ 78.400001n V_hig
+ 78.500000n V_hig
+ 78.500001n V_hig
+ 78.600000n V_hig
+ 78.600001n V_hig
+ 78.700000n V_hig
+ 78.700001n V_hig
+ 78.800000n V_hig
+ 78.800001n V_hig
+ 78.900000n V_hig
+ 78.900001n V_hig
+ 79.000000n V_hig
+ 79.000001n V_low
+ 79.100000n V_low
+ 79.100001n V_low
+ 79.200000n V_low
+ 79.200001n V_low
+ 79.300000n V_low
+ 79.300001n V_low
+ 79.400000n V_low
+ 79.400001n V_low
+ 79.500000n V_low
+ 79.500001n V_low
+ 79.600000n V_low
+ 79.600001n V_low
+ 79.700000n V_low
+ 79.700001n V_low
+ 79.800000n V_low
+ 79.800001n V_low
+ 79.900000n V_low
+ 79.900001n V_low
+ 80.000000n V_low
+ 80.000001n V_hig
+ 80.100000n V_hig
+ 80.100001n V_hig
+ 80.200000n V_hig
+ 80.200001n V_hig
+ 80.300000n V_hig
+ 80.300001n V_hig
+ 80.400000n V_hig
+ 80.400001n V_hig
+ 80.500000n V_hig
+ 80.500001n V_hig
+ 80.600000n V_hig
+ 80.600001n V_hig
+ 80.700000n V_hig
+ 80.700001n V_hig
+ 80.800000n V_hig
+ 80.800001n V_hig
+ 80.900000n V_hig
+ 80.900001n V_hig
+ 81.000000n V_hig
+ 81.000001n V_low
+ 81.100000n V_low
+ 81.100001n V_low
+ 81.200000n V_low
+ 81.200001n V_low
+ 81.300000n V_low
+ 81.300001n V_low
+ 81.400000n V_low
+ 81.400001n V_low
+ 81.500000n V_low
+ 81.500001n V_low
+ 81.600000n V_low
+ 81.600001n V_low
+ 81.700000n V_low
+ 81.700001n V_low
+ 81.800000n V_low
+ 81.800001n V_low
+ 81.900000n V_low
+ 81.900001n V_low
+ 82.000000n V_low
+ 82.000001n V_hig
+ 82.100000n V_hig
+ 82.100001n V_hig
+ 82.200000n V_hig
+ 82.200001n V_hig
+ 82.300000n V_hig
+ 82.300001n V_hig
+ 82.400000n V_hig
+ 82.400001n V_hig
+ 82.500000n V_hig
+ 82.500001n V_hig
+ 82.600000n V_hig
+ 82.600001n V_hig
+ 82.700000n V_hig
+ 82.700001n V_hig
+ 82.800000n V_hig
+ 82.800001n V_hig
+ 82.900000n V_hig
+ 82.900001n V_hig
+ 83.000000n V_hig
+ 83.000001n V_low
+ 83.100000n V_low
+ 83.100001n V_low
+ 83.200000n V_low
+ 83.200001n V_low
+ 83.300000n V_low
+ 83.300001n V_low
+ 83.400000n V_low
+ 83.400001n V_low
+ 83.500000n V_low
+ 83.500001n V_low
+ 83.600000n V_low
+ 83.600001n V_low
+ 83.700000n V_low
+ 83.700001n V_low
+ 83.800000n V_low
+ 83.800001n V_low
+ 83.900000n V_low
+ 83.900001n V_low
+ 84.000000n V_low
+ 84.000001n V_hig
+ 84.100000n V_hig
+ 84.100001n V_hig
+ 84.200000n V_hig
+ 84.200001n V_hig
+ 84.300000n V_hig
+ 84.300001n V_hig
+ 84.400000n V_hig
+ 84.400001n V_hig
+ 84.500000n V_hig
+ 84.500001n V_hig
+ 84.600000n V_hig
+ 84.600001n V_hig
+ 84.700000n V_hig
+ 84.700001n V_hig
+ 84.800000n V_hig
+ 84.800001n V_hig
+ 84.900000n V_hig
+ 84.900001n V_hig
+ 85.000000n V_hig
+ 85.000001n V_hig
+ 85.100000n V_hig
+ 85.100001n V_hig
+ 85.200000n V_hig
+ 85.200001n V_hig
+ 85.300000n V_hig
+ 85.300001n V_hig
+ 85.400000n V_hig
+ 85.400001n V_hig
+ 85.500000n V_hig
+ 85.500001n V_hig
+ 85.600000n V_hig
+ 85.600001n V_hig
+ 85.700000n V_hig
+ 85.700001n V_hig
+ 85.800000n V_hig
+ 85.800001n V_hig
+ 85.900000n V_hig
+ 85.900001n V_hig
+ 86.000000n V_hig
+ 86.000001n V_hig
+ 86.100000n V_hig
+ 86.100001n V_hig
+ 86.200000n V_hig
+ 86.200001n V_hig
+ 86.300000n V_hig
+ 86.300001n V_hig
+ 86.400000n V_hig
+ 86.400001n V_hig
+ 86.500000n V_hig
+ 86.500001n V_hig
+ 86.600000n V_hig
+ 86.600001n V_hig
+ 86.700000n V_hig
+ 86.700001n V_hig
+ 86.800000n V_hig
+ 86.800001n V_hig
+ 86.900000n V_hig
+ 86.900001n V_hig
+ 87.000000n V_hig
+ 87.000001n V_hig
+ 87.100000n V_hig
+ 87.100001n V_hig
+ 87.200000n V_hig
+ 87.200001n V_hig
+ 87.300000n V_hig
+ 87.300001n V_hig
+ 87.400000n V_hig
+ 87.400001n V_hig
+ 87.500000n V_hig
+ 87.500001n V_hig
+ 87.600000n V_hig
+ 87.600001n V_hig
+ 87.700000n V_hig
+ 87.700001n V_hig
+ 87.800000n V_hig
+ 87.800001n V_hig
+ 87.900000n V_hig
+ 87.900001n V_hig
+ 88.000000n V_hig
+ 88.000001n V_hig
+ 88.100000n V_hig
+ 88.100001n V_hig
+ 88.200000n V_hig
+ 88.200001n V_hig
+ 88.300000n V_hig
+ 88.300001n V_hig
+ 88.400000n V_hig
+ 88.400001n V_hig
+ 88.500000n V_hig
+ 88.500001n V_hig
+ 88.600000n V_hig
+ 88.600001n V_hig
+ 88.700000n V_hig
+ 88.700001n V_hig
+ 88.800000n V_hig
+ 88.800001n V_hig
+ 88.900000n V_hig
+ 88.900001n V_hig
+ 89.000000n V_hig
+ 89.000001n V_low
+ 89.100000n V_low
+ 89.100001n V_low
+ 89.200000n V_low
+ 89.200001n V_low
+ 89.300000n V_low
+ 89.300001n V_low
+ 89.400000n V_low
+ 89.400001n V_low
+ 89.500000n V_low
+ 89.500001n V_low
+ 89.600000n V_low
+ 89.600001n V_low
+ 89.700000n V_low
+ 89.700001n V_low
+ 89.800000n V_low
+ 89.800001n V_low
+ 89.900000n V_low
+ 89.900001n V_low
+ 90.000000n V_low
+ 90.000001n V_hig
+ 90.100000n V_hig
+ 90.100001n V_hig
+ 90.200000n V_hig
+ 90.200001n V_hig
+ 90.300000n V_hig
+ 90.300001n V_hig
+ 90.400000n V_hig
+ 90.400001n V_hig
+ 90.500000n V_hig
+ 90.500001n V_hig
+ 90.600000n V_hig
+ 90.600001n V_hig
+ 90.700000n V_hig
+ 90.700001n V_hig
+ 90.800000n V_hig
+ 90.800001n V_hig
+ 90.900000n V_hig
+ 90.900001n V_hig
+ 91.000000n V_hig
+ 91.000001n V_hig
+ 91.100000n V_hig
+ 91.100001n V_hig
+ 91.200000n V_hig
+ 91.200001n V_hig
+ 91.300000n V_hig
+ 91.300001n V_hig
+ 91.400000n V_hig
+ 91.400001n V_hig
+ 91.500000n V_hig
+ 91.500001n V_hig
+ 91.600000n V_hig
+ 91.600001n V_hig
+ 91.700000n V_hig
+ 91.700001n V_hig
+ 91.800000n V_hig
+ 91.800001n V_hig
+ 91.900000n V_hig
+ 91.900001n V_hig
+ 92.000000n V_hig
+ 92.000001n V_low
+ 92.100000n V_low
+ 92.100001n V_low
+ 92.200000n V_low
+ 92.200001n V_low
+ 92.300000n V_low
+ 92.300001n V_low
+ 92.400000n V_low
+ 92.400001n V_low
+ 92.500000n V_low
+ 92.500001n V_low
+ 92.600000n V_low
+ 92.600001n V_low
+ 92.700000n V_low
+ 92.700001n V_low
+ 92.800000n V_low
+ 92.800001n V_low
+ 92.900000n V_low
+ 92.900001n V_low
+ 93.000000n V_low
+ 93.000001n V_low
+ 93.100000n V_low
+ 93.100001n V_low
+ 93.200000n V_low
+ 93.200001n V_low
+ 93.300000n V_low
+ 93.300001n V_low
+ 93.400000n V_low
+ 93.400001n V_low
+ 93.500000n V_low
+ 93.500001n V_low
+ 93.600000n V_low
+ 93.600001n V_low
+ 93.700000n V_low
+ 93.700001n V_low
+ 93.800000n V_low
+ 93.800001n V_low
+ 93.900000n V_low
+ 93.900001n V_low
+ 94.000000n V_low
+ 94.000001n V_hig
+ 94.100000n V_hig
+ 94.100001n V_hig
+ 94.200000n V_hig
+ 94.200001n V_hig
+ 94.300000n V_hig
+ 94.300001n V_hig
+ 94.400000n V_hig
+ 94.400001n V_hig
+ 94.500000n V_hig
+ 94.500001n V_hig
+ 94.600000n V_hig
+ 94.600001n V_hig
+ 94.700000n V_hig
+ 94.700001n V_hig
+ 94.800000n V_hig
+ 94.800001n V_hig
+ 94.900000n V_hig
+ 94.900001n V_hig
+ 95.000000n V_hig
+ 95.000001n V_hig
+ 95.100000n V_hig
+ 95.100001n V_hig
+ 95.200000n V_hig
+ 95.200001n V_hig
+ 95.300000n V_hig
+ 95.300001n V_hig
+ 95.400000n V_hig
+ 95.400001n V_hig
+ 95.500000n V_hig
+ 95.500001n V_hig
+ 95.600000n V_hig
+ 95.600001n V_hig
+ 95.700000n V_hig
+ 95.700001n V_hig
+ 95.800000n V_hig
+ 95.800001n V_hig
+ 95.900000n V_hig
+ 95.900001n V_hig
+ 96.000000n V_hig
+ 96.000001n V_hig
+ 96.100000n V_hig
+ 96.100001n V_hig
+ 96.200000n V_hig
+ 96.200001n V_hig
+ 96.300000n V_hig
+ 96.300001n V_hig
+ 96.400000n V_hig
+ 96.400001n V_hig
+ 96.500000n V_hig
+ 96.500001n V_hig
+ 96.600000n V_hig
+ 96.600001n V_hig
+ 96.700000n V_hig
+ 96.700001n V_hig
+ 96.800000n V_hig
+ 96.800001n V_hig
+ 96.900000n V_hig
+ 96.900001n V_hig
+ 97.000000n V_hig
+ 97.000001n V_low
+ 97.100000n V_low
+ 97.100001n V_low
+ 97.200000n V_low
+ 97.200001n V_low
+ 97.300000n V_low
+ 97.300001n V_low
+ 97.400000n V_low
+ 97.400001n V_low
+ 97.500000n V_low
+ 97.500001n V_low
+ 97.600000n V_low
+ 97.600001n V_low
+ 97.700000n V_low
+ 97.700001n V_low
+ 97.800000n V_low
+ 97.800001n V_low
+ 97.900000n V_low
+ 97.900001n V_low
+ 98.000000n V_low
+ 98.000001n V_hig
+ 98.100000n V_hig
+ 98.100001n V_hig
+ 98.200000n V_hig
+ 98.200001n V_hig
+ 98.300000n V_hig
+ 98.300001n V_hig
+ 98.400000n V_hig
+ 98.400001n V_hig
+ 98.500000n V_hig
+ 98.500001n V_hig
+ 98.600000n V_hig
+ 98.600001n V_hig
+ 98.700000n V_hig
+ 98.700001n V_hig
+ 98.800000n V_hig
+ 98.800001n V_hig
+ 98.900000n V_hig
+ 98.900001n V_hig
+ 99.000000n V_hig
+ 99.000001n V_hig
+ 99.100000n V_hig
+ 99.100001n V_hig
+ 99.200000n V_hig
+ 99.200001n V_hig
+ 99.300000n V_hig
+ 99.300001n V_hig
+ 99.400000n V_hig
+ 99.400001n V_hig
+ 99.500000n V_hig
+ 99.500001n V_hig
+ 99.600000n V_hig
+ 99.600001n V_hig
+ 99.700000n V_hig
+ 99.700001n V_hig
+ 99.800000n V_hig
+ 99.800001n V_hig
+ 99.900000n V_hig
+ 99.900001n V_hig
+ 100.000000n V_hig
+ 100.000001n V_hig
+ 100.100000n V_hig
+ 100.100001n V_hig
+ 100.200000n V_hig
+ 100.200001n V_hig
+ 100.300000n V_hig
+ 100.300001n V_hig
+ 100.400000n V_hig
+ 100.400001n V_hig
+ 100.500000n V_hig
+ 100.500001n V_hig
+ 100.600000n V_hig
+ 100.600001n V_hig
+ 100.700000n V_hig
+ 100.700001n V_hig
+ 100.800000n V_hig
+ 100.800001n V_hig
+ 100.900000n V_hig
+ 100.900001n V_hig
+ 101.000000n V_hig
+ 101.000001n V_low
+ 101.100000n V_low
+ 101.100001n V_low
+ 101.200000n V_low
+ 101.200001n V_low
+ 101.300000n V_low
+ 101.300001n V_low
+ 101.400000n V_low
+ 101.400001n V_low
+ 101.500000n V_low
+ 101.500001n V_low
+ 101.600000n V_low
+ 101.600001n V_low
+ 101.700000n V_low
+ 101.700001n V_low
+ 101.800000n V_low
+ 101.800001n V_low
+ 101.900000n V_low
+ 101.900001n V_low
+ 102.000000n V_low
+ 102.000001n V_hig
+ 102.100000n V_hig
+ 102.100001n V_hig
+ 102.200000n V_hig
+ 102.200001n V_hig
+ 102.300000n V_hig
+ 102.300001n V_hig
+ 102.400000n V_hig
+ 102.400001n V_hig
+ 102.500000n V_hig
+ 102.500001n V_hig
+ 102.600000n V_hig
+ 102.600001n V_hig
+ 102.700000n V_hig
+ 102.700001n V_hig
+ 102.800000n V_hig
+ 102.800001n V_hig
+ 102.900000n V_hig
+ 102.900001n V_hig
+ 103.000000n V_hig
+ 103.000001n V_hig
+ 103.100000n V_hig
+ 103.100001n V_hig
+ 103.200000n V_hig
+ 103.200001n V_hig
+ 103.300000n V_hig
+ 103.300001n V_hig
+ 103.400000n V_hig
+ 103.400001n V_hig
+ 103.500000n V_hig
+ 103.500001n V_hig
+ 103.600000n V_hig
+ 103.600001n V_hig
+ 103.700000n V_hig
+ 103.700001n V_hig
+ 103.800000n V_hig
+ 103.800001n V_hig
+ 103.900000n V_hig
+ 103.900001n V_hig
+ 104.000000n V_hig
+ 104.000001n V_hig
+ 104.100000n V_hig
+ 104.100001n V_hig
+ 104.200000n V_hig
+ 104.200001n V_hig
+ 104.300000n V_hig
+ 104.300001n V_hig
+ 104.400000n V_hig
+ 104.400001n V_hig
+ 104.500000n V_hig
+ 104.500001n V_hig
+ 104.600000n V_hig
+ 104.600001n V_hig
+ 104.700000n V_hig
+ 104.700001n V_hig
+ 104.800000n V_hig
+ 104.800001n V_hig
+ 104.900000n V_hig
+ 104.900001n V_hig
+ 105.000000n V_hig
+ 105.000001n V_hig
+ 105.100000n V_hig
+ 105.100001n V_hig
+ 105.200000n V_hig
+ 105.200001n V_hig
+ 105.300000n V_hig
+ 105.300001n V_hig
+ 105.400000n V_hig
+ 105.400001n V_hig
+ 105.500000n V_hig
+ 105.500001n V_hig
+ 105.600000n V_hig
+ 105.600001n V_hig
+ 105.700000n V_hig
+ 105.700001n V_hig
+ 105.800000n V_hig
+ 105.800001n V_hig
+ 105.900000n V_hig
+ 105.900001n V_hig
+ 106.000000n V_hig
+ 106.000001n V_hig
+ 106.100000n V_hig
+ 106.100001n V_hig
+ 106.200000n V_hig
+ 106.200001n V_hig
+ 106.300000n V_hig
+ 106.300001n V_hig
+ 106.400000n V_hig
+ 106.400001n V_hig
+ 106.500000n V_hig
+ 106.500001n V_hig
+ 106.600000n V_hig
+ 106.600001n V_hig
+ 106.700000n V_hig
+ 106.700001n V_hig
+ 106.800000n V_hig
+ 106.800001n V_hig
+ 106.900000n V_hig
+ 106.900001n V_hig
+ 107.000000n V_hig
+ 107.000001n V_hig
+ 107.100000n V_hig
+ 107.100001n V_hig
+ 107.200000n V_hig
+ 107.200001n V_hig
+ 107.300000n V_hig
+ 107.300001n V_hig
+ 107.400000n V_hig
+ 107.400001n V_hig
+ 107.500000n V_hig
+ 107.500001n V_hig
+ 107.600000n V_hig
+ 107.600001n V_hig
+ 107.700000n V_hig
+ 107.700001n V_hig
+ 107.800000n V_hig
+ 107.800001n V_hig
+ 107.900000n V_hig
+ 107.900001n V_hig
+ 108.000000n V_hig
+ 108.000001n V_hig
+ 108.100000n V_hig
+ 108.100001n V_hig
+ 108.200000n V_hig
+ 108.200001n V_hig
+ 108.300000n V_hig
+ 108.300001n V_hig
+ 108.400000n V_hig
+ 108.400001n V_hig
+ 108.500000n V_hig
+ 108.500001n V_hig
+ 108.600000n V_hig
+ 108.600001n V_hig
+ 108.700000n V_hig
+ 108.700001n V_hig
+ 108.800000n V_hig
+ 108.800001n V_hig
+ 108.900000n V_hig
+ 108.900001n V_hig
+ 109.000000n V_hig
+ 109.000001n V_low
+ 109.100000n V_low
+ 109.100001n V_low
+ 109.200000n V_low
+ 109.200001n V_low
+ 109.300000n V_low
+ 109.300001n V_low
+ 109.400000n V_low
+ 109.400001n V_low
+ 109.500000n V_low
+ 109.500001n V_low
+ 109.600000n V_low
+ 109.600001n V_low
+ 109.700000n V_low
+ 109.700001n V_low
+ 109.800000n V_low
+ 109.800001n V_low
+ 109.900000n V_low
+ 109.900001n V_low
+ 110.000000n V_low
+ 110.000001n V_hig
+ 110.100000n V_hig
+ 110.100001n V_hig
+ 110.200000n V_hig
+ 110.200001n V_hig
+ 110.300000n V_hig
+ 110.300001n V_hig
+ 110.400000n V_hig
+ 110.400001n V_hig
+ 110.500000n V_hig
+ 110.500001n V_hig
+ 110.600000n V_hig
+ 110.600001n V_hig
+ 110.700000n V_hig
+ 110.700001n V_hig
+ 110.800000n V_hig
+ 110.800001n V_hig
+ 110.900000n V_hig
+ 110.900001n V_hig
+ 111.000000n V_hig
+ 111.000001n V_hig
+ 111.100000n V_hig
+ 111.100001n V_hig
+ 111.200000n V_hig
+ 111.200001n V_hig
+ 111.300000n V_hig
+ 111.300001n V_hig
+ 111.400000n V_hig
+ 111.400001n V_hig
+ 111.500000n V_hig
+ 111.500001n V_hig
+ 111.600000n V_hig
+ 111.600001n V_hig
+ 111.700000n V_hig
+ 111.700001n V_hig
+ 111.800000n V_hig
+ 111.800001n V_hig
+ 111.900000n V_hig
+ 111.900001n V_hig
+ 112.000000n V_hig
+ 112.000001n V_hig
+ 112.100000n V_hig
+ 112.100001n V_hig
+ 112.200000n V_hig
+ 112.200001n V_hig
+ 112.300000n V_hig
+ 112.300001n V_hig
+ 112.400000n V_hig
+ 112.400001n V_hig
+ 112.500000n V_hig
+ 112.500001n V_hig
+ 112.600000n V_hig
+ 112.600001n V_hig
+ 112.700000n V_hig
+ 112.700001n V_hig
+ 112.800000n V_hig
+ 112.800001n V_hig
+ 112.900000n V_hig
+ 112.900001n V_hig
+ 113.000000n V_hig
+ 113.000001n V_low
+ 113.100000n V_low
+ 113.100001n V_low
+ 113.200000n V_low
+ 113.200001n V_low
+ 113.300000n V_low
+ 113.300001n V_low
+ 113.400000n V_low
+ 113.400001n V_low
+ 113.500000n V_low
+ 113.500001n V_low
+ 113.600000n V_low
+ 113.600001n V_low
+ 113.700000n V_low
+ 113.700001n V_low
+ 113.800000n V_low
+ 113.800001n V_low
+ 113.900000n V_low
+ 113.900001n V_low
+ 114.000000n V_low
+ 114.000001n V_low
+ 114.100000n V_low
+ 114.100001n V_low
+ 114.200000n V_low
+ 114.200001n V_low
+ 114.300000n V_low
+ 114.300001n V_low
+ 114.400000n V_low
+ 114.400001n V_low
+ 114.500000n V_low
+ 114.500001n V_low
+ 114.600000n V_low
+ 114.600001n V_low
+ 114.700000n V_low
+ 114.700001n V_low
+ 114.800000n V_low
+ 114.800001n V_low
+ 114.900000n V_low
+ 114.900001n V_low
+ 115.000000n V_low
+ 115.000001n V_low
+ 115.100000n V_low
+ 115.100001n V_low
+ 115.200000n V_low
+ 115.200001n V_low
+ 115.300000n V_low
+ 115.300001n V_low
+ 115.400000n V_low
+ 115.400001n V_low
+ 115.500000n V_low
+ 115.500001n V_low
+ 115.600000n V_low
+ 115.600001n V_low
+ 115.700000n V_low
+ 115.700001n V_low
+ 115.800000n V_low
+ 115.800001n V_low
+ 115.900000n V_low
+ 115.900001n V_low
+ 116.000000n V_low
+ 116.000001n V_hig
+ 116.100000n V_hig
+ 116.100001n V_hig
+ 116.200000n V_hig
+ 116.200001n V_hig
+ 116.300000n V_hig
+ 116.300001n V_hig
+ 116.400000n V_hig
+ 116.400001n V_hig
+ 116.500000n V_hig
+ 116.500001n V_hig
+ 116.600000n V_hig
+ 116.600001n V_hig
+ 116.700000n V_hig
+ 116.700001n V_hig
+ 116.800000n V_hig
+ 116.800001n V_hig
+ 116.900000n V_hig
+ 116.900001n V_hig
+ 117.000000n V_hig
+ 117.000001n V_low
+ 117.100000n V_low
+ 117.100001n V_low
+ 117.200000n V_low
+ 117.200001n V_low
+ 117.300000n V_low
+ 117.300001n V_low
+ 117.400000n V_low
+ 117.400001n V_low
+ 117.500000n V_low
+ 117.500001n V_low
+ 117.600000n V_low
+ 117.600001n V_low
+ 117.700000n V_low
+ 117.700001n V_low
+ 117.800000n V_low
+ 117.800001n V_low
+ 117.900000n V_low
+ 117.900001n V_low
+ 118.000000n V_low
+ 118.000001n V_low
+ 118.100000n V_low
+ 118.100001n V_low
+ 118.200000n V_low
+ 118.200001n V_low
+ 118.300000n V_low
+ 118.300001n V_low
+ 118.400000n V_low
+ 118.400001n V_low
+ 118.500000n V_low
+ 118.500001n V_low
+ 118.600000n V_low
+ 118.600001n V_low
+ 118.700000n V_low
+ 118.700001n V_low
+ 118.800000n V_low
+ 118.800001n V_low
+ 118.900000n V_low
+ 118.900001n V_low
+ 119.000000n V_low
+ 119.000001n V_hig
+ 119.100000n V_hig
+ 119.100001n V_hig
+ 119.200000n V_hig
+ 119.200001n V_hig
+ 119.300000n V_hig
+ 119.300001n V_hig
+ 119.400000n V_hig
+ 119.400001n V_hig
+ 119.500000n V_hig
+ 119.500001n V_hig
+ 119.600000n V_hig
+ 119.600001n V_hig
+ 119.700000n V_hig
+ 119.700001n V_hig
+ 119.800000n V_hig
+ 119.800001n V_hig
+ 119.900000n V_hig
+ 119.900001n V_hig
+ 120.000000n V_hig
+ 120.000001n V_hig
+ 120.100000n V_hig
+ 120.100001n V_hig
+ 120.200000n V_hig
+ 120.200001n V_hig
+ 120.300000n V_hig
+ 120.300001n V_hig
+ 120.400000n V_hig
+ 120.400001n V_hig
+ 120.500000n V_hig
+ 120.500001n V_hig
+ 120.600000n V_hig
+ 120.600001n V_hig
+ 120.700000n V_hig
+ 120.700001n V_hig
+ 120.800000n V_hig
+ 120.800001n V_hig
+ 120.900000n V_hig
+ 120.900001n V_hig
+ 121.000000n V_hig
+ 121.000001n V_low
+ 121.100000n V_low
+ 121.100001n V_low
+ 121.200000n V_low
+ 121.200001n V_low
+ 121.300000n V_low
+ 121.300001n V_low
+ 121.400000n V_low
+ 121.400001n V_low
+ 121.500000n V_low
+ 121.500001n V_low
+ 121.600000n V_low
+ 121.600001n V_low
+ 121.700000n V_low
+ 121.700001n V_low
+ 121.800000n V_low
+ 121.800001n V_low
+ 121.900000n V_low
+ 121.900001n V_low
+ 122.000000n V_low
+ 122.000001n V_hig
+ 122.100000n V_hig
+ 122.100001n V_hig
+ 122.200000n V_hig
+ 122.200001n V_hig
+ 122.300000n V_hig
+ 122.300001n V_hig
+ 122.400000n V_hig
+ 122.400001n V_hig
+ 122.500000n V_hig
+ 122.500001n V_hig
+ 122.600000n V_hig
+ 122.600001n V_hig
+ 122.700000n V_hig
+ 122.700001n V_hig
+ 122.800000n V_hig
+ 122.800001n V_hig
+ 122.900000n V_hig
+ 122.900001n V_hig
+ 123.000000n V_hig
+ 123.000001n V_low
+ 123.100000n V_low
+ 123.100001n V_low
+ 123.200000n V_low
+ 123.200001n V_low
+ 123.300000n V_low
+ 123.300001n V_low
+ 123.400000n V_low
+ 123.400001n V_low
+ 123.500000n V_low
+ 123.500001n V_low
+ 123.600000n V_low
+ 123.600001n V_low
+ 123.700000n V_low
+ 123.700001n V_low
+ 123.800000n V_low
+ 123.800001n V_low
+ 123.900000n V_low
+ 123.900001n V_low
+ 124.000000n V_low
+ 124.000001n V_low
+ 124.100000n V_low
+ 124.100001n V_low
+ 124.200000n V_low
+ 124.200001n V_low
+ 124.300000n V_low
+ 124.300001n V_low
+ 124.400000n V_low
+ 124.400001n V_low
+ 124.500000n V_low
+ 124.500001n V_low
+ 124.600000n V_low
+ 124.600001n V_low
+ 124.700000n V_low
+ 124.700001n V_low
+ 124.800000n V_low
+ 124.800001n V_low
+ 124.900000n V_low
+ 124.900001n V_low
+ 125.000000n V_low
+ 125.000001n V_low
+ 125.100000n V_low
+ 125.100001n V_low
+ 125.200000n V_low
+ 125.200001n V_low
+ 125.300000n V_low
+ 125.300001n V_low
+ 125.400000n V_low
+ 125.400001n V_low
+ 125.500000n V_low
+ 125.500001n V_low
+ 125.600000n V_low
+ 125.600001n V_low
+ 125.700000n V_low
+ 125.700001n V_low
+ 125.800000n V_low
+ 125.800001n V_low
+ 125.900000n V_low
+ 125.900001n V_low
+ 126.000000n V_low
+ 126.000001n V_hig
+ 126.100000n V_hig
+ 126.100001n V_hig
+ 126.200000n V_hig
+ 126.200001n V_hig
+ 126.300000n V_hig
+ 126.300001n V_hig
+ 126.400000n V_hig
+ 126.400001n V_hig
+ 126.500000n V_hig
+ 126.500001n V_hig
+ 126.600000n V_hig
+ 126.600001n V_hig
+ 126.700000n V_hig
+ 126.700001n V_hig
+ 126.800000n V_hig
+ 126.800001n V_hig
+ 126.900000n V_hig
+ 126.900001n V_hig
+ 127.000000n V_hig
+ 127.000001n V_low
+ 127.100000n V_low
+ 127.100001n V_low
+ 127.200000n V_low
+ 127.200001n V_low
+ 127.300000n V_low
+ 127.300001n V_low
+ 127.400000n V_low
+ 127.400001n V_low
+ 127.500000n V_low
+ 127.500001n V_low
+ 127.600000n V_low
+ 127.600001n V_low
+ 127.700000n V_low
+ 127.700001n V_low
+ 127.800000n V_low
+ 127.800001n V_low
+ 127.900000n V_low
+ 127.900001n V_low
+ 128.000000n V_low
+ 128.000001n V_low
+ 128.100000n V_low
+ 128.100001n V_low
+ 128.200000n V_low
+ 128.200001n V_low
+ 128.300000n V_low
+ 128.300001n V_low
+ 128.400000n V_low
+ 128.400001n V_low
+ 128.500000n V_low
+ 128.500001n V_low
+ 128.600000n V_low
+ 128.600001n V_low
+ 128.700000n V_low
+ 128.700001n V_low
+ 128.800000n V_low
+ 128.800001n V_low
+ 128.900000n V_low
+ 128.900001n V_low
+ 129.000000n V_low
+ 129.000001n V_low
+ 129.100000n V_low
+ 129.100001n V_low
+ 129.200000n V_low
+ 129.200001n V_low
+ 129.300000n V_low
+ 129.300001n V_low
+ 129.400000n V_low
+ 129.400001n V_low
+ 129.500000n V_low
+ 129.500001n V_low
+ 129.600000n V_low
+ 129.600001n V_low
+ 129.700000n V_low
+ 129.700001n V_low
+ 129.800000n V_low
+ 129.800001n V_low
+ 129.900000n V_low
+ 129.900001n V_low
+ 130.000000n V_low
+ 130.000001n V_low
+ 130.100000n V_low
+ 130.100001n V_low
+ 130.200000n V_low
+ 130.200001n V_low
+ 130.300000n V_low
+ 130.300001n V_low
+ 130.400000n V_low
+ 130.400001n V_low
+ 130.500000n V_low
+ 130.500001n V_low
+ 130.600000n V_low
+ 130.600001n V_low
+ 130.700000n V_low
+ 130.700001n V_low
+ 130.800000n V_low
+ 130.800001n V_low
+ 130.900000n V_low
+ 130.900001n V_low
+ 131.000000n V_low
+ 131.000001n V_low
+ 131.100000n V_low
+ 131.100001n V_low
+ 131.200000n V_low
+ 131.200001n V_low
+ 131.300000n V_low
+ 131.300001n V_low
+ 131.400000n V_low
+ 131.400001n V_low
+ 131.500000n V_low
+ 131.500001n V_low
+ 131.600000n V_low
+ 131.600001n V_low
+ 131.700000n V_low
+ 131.700001n V_low
+ 131.800000n V_low
+ 131.800001n V_low
+ 131.900000n V_low
+ 131.900001n V_low
+ 132.000000n V_low
+ 132.000001n V_low
+ 132.100000n V_low
+ 132.100001n V_low
+ 132.200000n V_low
+ 132.200001n V_low
+ 132.300000n V_low
+ 132.300001n V_low
+ 132.400000n V_low
+ 132.400001n V_low
+ 132.500000n V_low
+ 132.500001n V_low
+ 132.600000n V_low
+ 132.600001n V_low
+ 132.700000n V_low
+ 132.700001n V_low
+ 132.800000n V_low
+ 132.800001n V_low
+ 132.900000n V_low
+ 132.900001n V_low
+ 133.000000n V_low
+ 133.000001n V_low
+ 133.100000n V_low
+ 133.100001n V_low
+ 133.200000n V_low
+ 133.200001n V_low
+ 133.300000n V_low
+ 133.300001n V_low
+ 133.400000n V_low
+ 133.400001n V_low
+ 133.500000n V_low
+ 133.500001n V_low
+ 133.600000n V_low
+ 133.600001n V_low
+ 133.700000n V_low
+ 133.700001n V_low
+ 133.800000n V_low
+ 133.800001n V_low
+ 133.900000n V_low
+ 133.900001n V_low
+ 134.000000n V_low
+ 134.000001n V_hig
+ 134.100000n V_hig
+ 134.100001n V_hig
+ 134.200000n V_hig
+ 134.200001n V_hig
+ 134.300000n V_hig
+ 134.300001n V_hig
+ 134.400000n V_hig
+ 134.400001n V_hig
+ 134.500000n V_hig
+ 134.500001n V_hig
+ 134.600000n V_hig
+ 134.600001n V_hig
+ 134.700000n V_hig
+ 134.700001n V_hig
+ 134.800000n V_hig
+ 134.800001n V_hig
+ 134.900000n V_hig
+ 134.900001n V_hig
+ 135.000000n V_hig
+ 135.000001n V_low
+ 135.100000n V_low
+ 135.100001n V_low
+ 135.200000n V_low
+ 135.200001n V_low
+ 135.300000n V_low
+ 135.300001n V_low
+ 135.400000n V_low
+ 135.400001n V_low
+ 135.500000n V_low
+ 135.500001n V_low
+ 135.600000n V_low
+ 135.600001n V_low
+ 135.700000n V_low
+ 135.700001n V_low
+ 135.800000n V_low
+ 135.800001n V_low
+ 135.900000n V_low
+ 135.900001n V_low
+ 136.000000n V_low
+ 136.000001n V_hig
+ 136.100000n V_hig
+ 136.100001n V_hig
+ 136.200000n V_hig
+ 136.200001n V_hig
+ 136.300000n V_hig
+ 136.300001n V_hig
+ 136.400000n V_hig
+ 136.400001n V_hig
+ 136.500000n V_hig
+ 136.500001n V_hig
+ 136.600000n V_hig
+ 136.600001n V_hig
+ 136.700000n V_hig
+ 136.700001n V_hig
+ 136.800000n V_hig
+ 136.800001n V_hig
+ 136.900000n V_hig
+ 136.900001n V_hig
+ 137.000000n V_hig
+ 137.000001n V_hig
+ 137.100000n V_hig
+ 137.100001n V_hig
+ 137.200000n V_hig
+ 137.200001n V_hig
+ 137.300000n V_hig
+ 137.300001n V_hig
+ 137.400000n V_hig
+ 137.400001n V_hig
+ 137.500000n V_hig
+ 137.500001n V_hig
+ 137.600000n V_hig
+ 137.600001n V_hig
+ 137.700000n V_hig
+ 137.700001n V_hig
+ 137.800000n V_hig
+ 137.800001n V_hig
+ 137.900000n V_hig
+ 137.900001n V_hig
+ 138.000000n V_hig
+ 138.000001n V_low
+ 138.100000n V_low
+ 138.100001n V_low
+ 138.200000n V_low
+ 138.200001n V_low
+ 138.300000n V_low
+ 138.300001n V_low
+ 138.400000n V_low
+ 138.400001n V_low
+ 138.500000n V_low
+ 138.500001n V_low
+ 138.600000n V_low
+ 138.600001n V_low
+ 138.700000n V_low
+ 138.700001n V_low
+ 138.800000n V_low
+ 138.800001n V_low
+ 138.900000n V_low
+ 138.900001n V_low
+ 139.000000n V_low
+ 139.000001n V_low
+ 139.100000n V_low
+ 139.100001n V_low
+ 139.200000n V_low
+ 139.200001n V_low
+ 139.300000n V_low
+ 139.300001n V_low
+ 139.400000n V_low
+ 139.400001n V_low
+ 139.500000n V_low
+ 139.500001n V_low
+ 139.600000n V_low
+ 139.600001n V_low
+ 139.700000n V_low
+ 139.700001n V_low
+ 139.800000n V_low
+ 139.800001n V_low
+ 139.900000n V_low
+ 139.900001n V_low
+ 140.000000n V_low
+ 140.000001n V_low
+ 140.100000n V_low
+ 140.100001n V_low
+ 140.200000n V_low
+ 140.200001n V_low
+ 140.300000n V_low
+ 140.300001n V_low
+ 140.400000n V_low
+ 140.400001n V_low
+ 140.500000n V_low
+ 140.500001n V_low
+ 140.600000n V_low
+ 140.600001n V_low
+ 140.700000n V_low
+ 140.700001n V_low
+ 140.800000n V_low
+ 140.800001n V_low
+ 140.900000n V_low
+ 140.900001n V_low
+ 141.000000n V_low
+ 141.000001n V_low
+ 141.100000n V_low
+ 141.100001n V_low
+ 141.200000n V_low
+ 141.200001n V_low
+ 141.300000n V_low
+ 141.300001n V_low
+ 141.400000n V_low
+ 141.400001n V_low
+ 141.500000n V_low
+ 141.500001n V_low
+ 141.600000n V_low
+ 141.600001n V_low
+ 141.700000n V_low
+ 141.700001n V_low
+ 141.800000n V_low
+ 141.800001n V_low
+ 141.900000n V_low
+ 141.900001n V_low
+ 142.000000n V_low
+ 142.000001n V_low
+ 142.100000n V_low
+ 142.100001n V_low
+ 142.200000n V_low
+ 142.200001n V_low
+ 142.300000n V_low
+ 142.300001n V_low
+ 142.400000n V_low
+ 142.400001n V_low
+ 142.500000n V_low
+ 142.500001n V_low
+ 142.600000n V_low
+ 142.600001n V_low
+ 142.700000n V_low
+ 142.700001n V_low
+ 142.800000n V_low
+ 142.800001n V_low
+ 142.900000n V_low
+ 142.900001n V_low
+ 143.000000n V_low
+ 143.000001n V_hig
+ 143.100000n V_hig
+ 143.100001n V_hig
+ 143.200000n V_hig
+ 143.200001n V_hig
+ 143.300000n V_hig
+ 143.300001n V_hig
+ 143.400000n V_hig
+ 143.400001n V_hig
+ 143.500000n V_hig
+ 143.500001n V_hig
+ 143.600000n V_hig
+ 143.600001n V_hig
+ 143.700000n V_hig
+ 143.700001n V_hig
+ 143.800000n V_hig
+ 143.800001n V_hig
+ 143.900000n V_hig
+ 143.900001n V_hig
+ 144.000000n V_hig
+ 144.000001n V_low
+ 144.100000n V_low
+ 144.100001n V_low
+ 144.200000n V_low
+ 144.200001n V_low
+ 144.300000n V_low
+ 144.300001n V_low
+ 144.400000n V_low
+ 144.400001n V_low
+ 144.500000n V_low
+ 144.500001n V_low
+ 144.600000n V_low
+ 144.600001n V_low
+ 144.700000n V_low
+ 144.700001n V_low
+ 144.800000n V_low
+ 144.800001n V_low
+ 144.900000n V_low
+ 144.900001n V_low
+ 145.000000n V_low
+ 145.000001n V_hig
+ 145.100000n V_hig
+ 145.100001n V_hig
+ 145.200000n V_hig
+ 145.200001n V_hig
+ 145.300000n V_hig
+ 145.300001n V_hig
+ 145.400000n V_hig
+ 145.400001n V_hig
+ 145.500000n V_hig
+ 145.500001n V_hig
+ 145.600000n V_hig
+ 145.600001n V_hig
+ 145.700000n V_hig
+ 145.700001n V_hig
+ 145.800000n V_hig
+ 145.800001n V_hig
+ 145.900000n V_hig
+ 145.900001n V_hig
+ 146.000000n V_hig
+ 146.000001n V_low
+ 146.100000n V_low
+ 146.100001n V_low
+ 146.200000n V_low
+ 146.200001n V_low
+ 146.300000n V_low
+ 146.300001n V_low
+ 146.400000n V_low
+ 146.400001n V_low
+ 146.500000n V_low
+ 146.500001n V_low
+ 146.600000n V_low
+ 146.600001n V_low
+ 146.700000n V_low
+ 146.700001n V_low
+ 146.800000n V_low
+ 146.800001n V_low
+ 146.900000n V_low
+ 146.900001n V_low
+ 147.000000n V_low
+ 147.000001n V_hig
+ 147.100000n V_hig
+ 147.100001n V_hig
+ 147.200000n V_hig
+ 147.200001n V_hig
+ 147.300000n V_hig
+ 147.300001n V_hig
+ 147.400000n V_hig
+ 147.400001n V_hig
+ 147.500000n V_hig
+ 147.500001n V_hig
+ 147.600000n V_hig
+ 147.600001n V_hig
+ 147.700000n V_hig
+ 147.700001n V_hig
+ 147.800000n V_hig
+ 147.800001n V_hig
+ 147.900000n V_hig
+ 147.900001n V_hig
+ 148.000000n V_hig
+ 148.000001n V_hig
+ 148.100000n V_hig
+ 148.100001n V_hig
+ 148.200000n V_hig
+ 148.200001n V_hig
+ 148.300000n V_hig
+ 148.300001n V_hig
+ 148.400000n V_hig
+ 148.400001n V_hig
+ 148.500000n V_hig
+ 148.500001n V_hig
+ 148.600000n V_hig
+ 148.600001n V_hig
+ 148.700000n V_hig
+ 148.700001n V_hig
+ 148.800000n V_hig
+ 148.800001n V_hig
+ 148.900000n V_hig
+ 148.900001n V_hig
+ 149.000000n V_hig
+ 149.000001n V_hig
+ 149.100000n V_hig
+ 149.100001n V_hig
+ 149.200000n V_hig
+ 149.200001n V_hig
+ 149.300000n V_hig
+ 149.300001n V_hig
+ 149.400000n V_hig
+ 149.400001n V_hig
+ 149.500000n V_hig
+ 149.500001n V_hig
+ 149.600000n V_hig
+ 149.600001n V_hig
+ 149.700000n V_hig
+ 149.700001n V_hig
+ 149.800000n V_hig
+ 149.800001n V_hig
+ 149.900000n V_hig
+ 149.900001n V_hig
+ 150.000000n V_hig
+ 150.000001n V_low
+ 150.100000n V_low
+ 150.100001n V_low
+ 150.200000n V_low
+ 150.200001n V_low
+ 150.300000n V_low
+ 150.300001n V_low
+ 150.400000n V_low
+ 150.400001n V_low
+ 150.500000n V_low
+ 150.500001n V_low
+ 150.600000n V_low
+ 150.600001n V_low
+ 150.700000n V_low
+ 150.700001n V_low
+ 150.800000n V_low
+ 150.800001n V_low
+ 150.900000n V_low
+ 150.900001n V_low
+ 151.000000n V_low
+ 151.000001n V_low
+ 151.100000n V_low
+ 151.100001n V_low
+ 151.200000n V_low
+ 151.200001n V_low
+ 151.300000n V_low
+ 151.300001n V_low
+ 151.400000n V_low
+ 151.400001n V_low
+ 151.500000n V_low
+ 151.500001n V_low
+ 151.600000n V_low
+ 151.600001n V_low
+ 151.700000n V_low
+ 151.700001n V_low
+ 151.800000n V_low
+ 151.800001n V_low
+ 151.900000n V_low
+ 151.900001n V_low
+ 152.000000n V_low
+ 152.000001n V_hig
+ 152.100000n V_hig
+ 152.100001n V_hig
+ 152.200000n V_hig
+ 152.200001n V_hig
+ 152.300000n V_hig
+ 152.300001n V_hig
+ 152.400000n V_hig
+ 152.400001n V_hig
+ 152.500000n V_hig
+ 152.500001n V_hig
+ 152.600000n V_hig
+ 152.600001n V_hig
+ 152.700000n V_hig
+ 152.700001n V_hig
+ 152.800000n V_hig
+ 152.800001n V_hig
+ 152.900000n V_hig
+ 152.900001n V_hig
+ 153.000000n V_hig
+ 153.000001n V_low
+ 153.100000n V_low
+ 153.100001n V_low
+ 153.200000n V_low
+ 153.200001n V_low
+ 153.300000n V_low
+ 153.300001n V_low
+ 153.400000n V_low
+ 153.400001n V_low
+ 153.500000n V_low
+ 153.500001n V_low
+ 153.600000n V_low
+ 153.600001n V_low
+ 153.700000n V_low
+ 153.700001n V_low
+ 153.800000n V_low
+ 153.800001n V_low
+ 153.900000n V_low
+ 153.900001n V_low
+ 154.000000n V_low
+ 154.000001n V_low
+ 154.100000n V_low
+ 154.100001n V_low
+ 154.200000n V_low
+ 154.200001n V_low
+ 154.300000n V_low
+ 154.300001n V_low
+ 154.400000n V_low
+ 154.400001n V_low
+ 154.500000n V_low
+ 154.500001n V_low
+ 154.600000n V_low
+ 154.600001n V_low
+ 154.700000n V_low
+ 154.700001n V_low
+ 154.800000n V_low
+ 154.800001n V_low
+ 154.900000n V_low
+ 154.900001n V_low
+ 155.000000n V_low
+ 155.000001n V_low
+ 155.100000n V_low
+ 155.100001n V_low
+ 155.200000n V_low
+ 155.200001n V_low
+ 155.300000n V_low
+ 155.300001n V_low
+ 155.400000n V_low
+ 155.400001n V_low
+ 155.500000n V_low
+ 155.500001n V_low
+ 155.600000n V_low
+ 155.600001n V_low
+ 155.700000n V_low
+ 155.700001n V_low
+ 155.800000n V_low
+ 155.800001n V_low
+ 155.900000n V_low
+ 155.900001n V_low
+ 156.000000n V_low
+ 156.000001n V_low
+ 156.100000n V_low
+ 156.100001n V_low
+ 156.200000n V_low
+ 156.200001n V_low
+ 156.300000n V_low
+ 156.300001n V_low
+ 156.400000n V_low
+ 156.400001n V_low
+ 156.500000n V_low
+ 156.500001n V_low
+ 156.600000n V_low
+ 156.600001n V_low
+ 156.700000n V_low
+ 156.700001n V_low
+ 156.800000n V_low
+ 156.800001n V_low
+ 156.900000n V_low
+ 156.900001n V_low
+ 157.000000n V_low
+ 157.000001n V_low
+ 157.100000n V_low
+ 157.100001n V_low
+ 157.200000n V_low
+ 157.200001n V_low
+ 157.300000n V_low
+ 157.300001n V_low
+ 157.400000n V_low
+ 157.400001n V_low
+ 157.500000n V_low
+ 157.500001n V_low
+ 157.600000n V_low
+ 157.600001n V_low
+ 157.700000n V_low
+ 157.700001n V_low
+ 157.800000n V_low
+ 157.800001n V_low
+ 157.900000n V_low
+ 157.900001n V_low
+ 158.000000n V_low
+ 158.000001n V_low
+ 158.100000n V_low
+ 158.100001n V_low
+ 158.200000n V_low
+ 158.200001n V_low
+ 158.300000n V_low
+ 158.300001n V_low
+ 158.400000n V_low
+ 158.400001n V_low
+ 158.500000n V_low
+ 158.500001n V_low
+ 158.600000n V_low
+ 158.600001n V_low
+ 158.700000n V_low
+ 158.700001n V_low
+ 158.800000n V_low
+ 158.800001n V_low
+ 158.900000n V_low
+ 158.900001n V_low
+ 159.000000n V_low
+ 159.000001n V_hig
+ 159.100000n V_hig
+ 159.100001n V_hig
+ 159.200000n V_hig
+ 159.200001n V_hig
+ 159.300000n V_hig
+ 159.300001n V_hig
+ 159.400000n V_hig
+ 159.400001n V_hig
+ 159.500000n V_hig
+ 159.500001n V_hig
+ 159.600000n V_hig
+ 159.600001n V_hig
+ 159.700000n V_hig
+ 159.700001n V_hig
+ 159.800000n V_hig
+ 159.800001n V_hig
+ 159.900000n V_hig
+ 159.900001n V_hig
+ 160.000000n V_hig
+ 160.000001n V_hig
+ 160.100000n V_hig
+ 160.100001n V_hig
+ 160.200000n V_hig
+ 160.200001n V_hig
+ 160.300000n V_hig
+ 160.300001n V_hig
+ 160.400000n V_hig
+ 160.400001n V_hig
+ 160.500000n V_hig
+ 160.500001n V_hig
+ 160.600000n V_hig
+ 160.600001n V_hig
+ 160.700000n V_hig
+ 160.700001n V_hig
+ 160.800000n V_hig
+ 160.800001n V_hig
+ 160.900000n V_hig
+ 160.900001n V_hig
+ 161.000000n V_hig
+ 161.000001n V_low
+ 161.100000n V_low
+ 161.100001n V_low
+ 161.200000n V_low
+ 161.200001n V_low
+ 161.300000n V_low
+ 161.300001n V_low
+ 161.400000n V_low
+ 161.400001n V_low
+ 161.500000n V_low
+ 161.500001n V_low
+ 161.600000n V_low
+ 161.600001n V_low
+ 161.700000n V_low
+ 161.700001n V_low
+ 161.800000n V_low
+ 161.800001n V_low
+ 161.900000n V_low
+ 161.900001n V_low
+ 162.000000n V_low
+ 162.000001n V_low
+ 162.100000n V_low
+ 162.100001n V_low
+ 162.200000n V_low
+ 162.200001n V_low
+ 162.300000n V_low
+ 162.300001n V_low
+ 162.400000n V_low
+ 162.400001n V_low
+ 162.500000n V_low
+ 162.500001n V_low
+ 162.600000n V_low
+ 162.600001n V_low
+ 162.700000n V_low
+ 162.700001n V_low
+ 162.800000n V_low
+ 162.800001n V_low
+ 162.900000n V_low
+ 162.900001n V_low
+ 163.000000n V_low
+ 163.000001n V_hig
+ 163.100000n V_hig
+ 163.100001n V_hig
+ 163.200000n V_hig
+ 163.200001n V_hig
+ 163.300000n V_hig
+ 163.300001n V_hig
+ 163.400000n V_hig
+ 163.400001n V_hig
+ 163.500000n V_hig
+ 163.500001n V_hig
+ 163.600000n V_hig
+ 163.600001n V_hig
+ 163.700000n V_hig
+ 163.700001n V_hig
+ 163.800000n V_hig
+ 163.800001n V_hig
+ 163.900000n V_hig
+ 163.900001n V_hig
+ 164.000000n V_hig
+ 164.000001n V_low
+ 164.100000n V_low
+ 164.100001n V_low
+ 164.200000n V_low
+ 164.200001n V_low
+ 164.300000n V_low
+ 164.300001n V_low
+ 164.400000n V_low
+ 164.400001n V_low
+ 164.500000n V_low
+ 164.500001n V_low
+ 164.600000n V_low
+ 164.600001n V_low
+ 164.700000n V_low
+ 164.700001n V_low
+ 164.800000n V_low
+ 164.800001n V_low
+ 164.900000n V_low
+ 164.900001n V_low
+ 165.000000n V_low
+ 165.000001n V_low
+ 165.100000n V_low
+ 165.100001n V_low
+ 165.200000n V_low
+ 165.200001n V_low
+ 165.300000n V_low
+ 165.300001n V_low
+ 165.400000n V_low
+ 165.400001n V_low
+ 165.500000n V_low
+ 165.500001n V_low
+ 165.600000n V_low
+ 165.600001n V_low
+ 165.700000n V_low
+ 165.700001n V_low
+ 165.800000n V_low
+ 165.800001n V_low
+ 165.900000n V_low
+ 165.900001n V_low
+ 166.000000n V_low
+ 166.000001n V_hig
+ 166.100000n V_hig
+ 166.100001n V_hig
+ 166.200000n V_hig
+ 166.200001n V_hig
+ 166.300000n V_hig
+ 166.300001n V_hig
+ 166.400000n V_hig
+ 166.400001n V_hig
+ 166.500000n V_hig
+ 166.500001n V_hig
+ 166.600000n V_hig
+ 166.600001n V_hig
+ 166.700000n V_hig
+ 166.700001n V_hig
+ 166.800000n V_hig
+ 166.800001n V_hig
+ 166.900000n V_hig
+ 166.900001n V_hig
+ 167.000000n V_hig
+ 167.000001n V_low
+ 167.100000n V_low
+ 167.100001n V_low
+ 167.200000n V_low
+ 167.200001n V_low
+ 167.300000n V_low
+ 167.300001n V_low
+ 167.400000n V_low
+ 167.400001n V_low
+ 167.500000n V_low
+ 167.500001n V_low
+ 167.600000n V_low
+ 167.600001n V_low
+ 167.700000n V_low
+ 167.700001n V_low
+ 167.800000n V_low
+ 167.800001n V_low
+ 167.900000n V_low
+ 167.900001n V_low
+ 168.000000n V_low
+ 168.000001n V_hig
+ 168.100000n V_hig
+ 168.100001n V_hig
+ 168.200000n V_hig
+ 168.200001n V_hig
+ 168.300000n V_hig
+ 168.300001n V_hig
+ 168.400000n V_hig
+ 168.400001n V_hig
+ 168.500000n V_hig
+ 168.500001n V_hig
+ 168.600000n V_hig
+ 168.600001n V_hig
+ 168.700000n V_hig
+ 168.700001n V_hig
+ 168.800000n V_hig
+ 168.800001n V_hig
+ 168.900000n V_hig
+ 168.900001n V_hig
+ 169.000000n V_hig
+ 169.000001n V_hig
+ 169.100000n V_hig
+ 169.100001n V_hig
+ 169.200000n V_hig
+ 169.200001n V_hig
+ 169.300000n V_hig
+ 169.300001n V_hig
+ 169.400000n V_hig
+ 169.400001n V_hig
+ 169.500000n V_hig
+ 169.500001n V_hig
+ 169.600000n V_hig
+ 169.600001n V_hig
+ 169.700000n V_hig
+ 169.700001n V_hig
+ 169.800000n V_hig
+ 169.800001n V_hig
+ 169.900000n V_hig
+ 169.900001n V_hig
+ 170.000000n V_hig
+ 170.000001n V_hig
+ 170.100000n V_hig
+ 170.100001n V_hig
+ 170.200000n V_hig
+ 170.200001n V_hig
+ 170.300000n V_hig
+ 170.300001n V_hig
+ 170.400000n V_hig
+ 170.400001n V_hig
+ 170.500000n V_hig
+ 170.500001n V_hig
+ 170.600000n V_hig
+ 170.600001n V_hig
+ 170.700000n V_hig
+ 170.700001n V_hig
+ 170.800000n V_hig
+ 170.800001n V_hig
+ 170.900000n V_hig
+ 170.900001n V_hig
+ 171.000000n V_hig
+ 171.000001n V_low
+ 171.100000n V_low
+ 171.100001n V_low
+ 171.200000n V_low
+ 171.200001n V_low
+ 171.300000n V_low
+ 171.300001n V_low
+ 171.400000n V_low
+ 171.400001n V_low
+ 171.500000n V_low
+ 171.500001n V_low
+ 171.600000n V_low
+ 171.600001n V_low
+ 171.700000n V_low
+ 171.700001n V_low
+ 171.800000n V_low
+ 171.800001n V_low
+ 171.900000n V_low
+ 171.900001n V_low
+ 172.000000n V_low
+ 172.000001n V_low
+ 172.100000n V_low
+ 172.100001n V_low
+ 172.200000n V_low
+ 172.200001n V_low
+ 172.300000n V_low
+ 172.300001n V_low
+ 172.400000n V_low
+ 172.400001n V_low
+ 172.500000n V_low
+ 172.500001n V_low
+ 172.600000n V_low
+ 172.600001n V_low
+ 172.700000n V_low
+ 172.700001n V_low
+ 172.800000n V_low
+ 172.800001n V_low
+ 172.900000n V_low
+ 172.900001n V_low
+ 173.000000n V_low
+ 173.000001n V_hig
+ 173.100000n V_hig
+ 173.100001n V_hig
+ 173.200000n V_hig
+ 173.200001n V_hig
+ 173.300000n V_hig
+ 173.300001n V_hig
+ 173.400000n V_hig
+ 173.400001n V_hig
+ 173.500000n V_hig
+ 173.500001n V_hig
+ 173.600000n V_hig
+ 173.600001n V_hig
+ 173.700000n V_hig
+ 173.700001n V_hig
+ 173.800000n V_hig
+ 173.800001n V_hig
+ 173.900000n V_hig
+ 173.900001n V_hig
+ 174.000000n V_hig
+ 174.000001n V_low
+ 174.100000n V_low
+ 174.100001n V_low
+ 174.200000n V_low
+ 174.200001n V_low
+ 174.300000n V_low
+ 174.300001n V_low
+ 174.400000n V_low
+ 174.400001n V_low
+ 174.500000n V_low
+ 174.500001n V_low
+ 174.600000n V_low
+ 174.600001n V_low
+ 174.700000n V_low
+ 174.700001n V_low
+ 174.800000n V_low
+ 174.800001n V_low
+ 174.900000n V_low
+ 174.900001n V_low
+ 175.000000n V_low
+ 175.000001n V_low
+ 175.100000n V_low
+ 175.100001n V_low
+ 175.200000n V_low
+ 175.200001n V_low
+ 175.300000n V_low
+ 175.300001n V_low
+ 175.400000n V_low
+ 175.400001n V_low
+ 175.500000n V_low
+ 175.500001n V_low
+ 175.600000n V_low
+ 175.600001n V_low
+ 175.700000n V_low
+ 175.700001n V_low
+ 175.800000n V_low
+ 175.800001n V_low
+ 175.900000n V_low
+ 175.900001n V_low
+ 176.000000n V_low
+ 176.000001n V_hig
+ 176.100000n V_hig
+ 176.100001n V_hig
+ 176.200000n V_hig
+ 176.200001n V_hig
+ 176.300000n V_hig
+ 176.300001n V_hig
+ 176.400000n V_hig
+ 176.400001n V_hig
+ 176.500000n V_hig
+ 176.500001n V_hig
+ 176.600000n V_hig
+ 176.600001n V_hig
+ 176.700000n V_hig
+ 176.700001n V_hig
+ 176.800000n V_hig
+ 176.800001n V_hig
+ 176.900000n V_hig
+ 176.900001n V_hig
+ 177.000000n V_hig
+ 177.000001n V_low
+ 177.100000n V_low
+ 177.100001n V_low
+ 177.200000n V_low
+ 177.200001n V_low
+ 177.300000n V_low
+ 177.300001n V_low
+ 177.400000n V_low
+ 177.400001n V_low
+ 177.500000n V_low
+ 177.500001n V_low
+ 177.600000n V_low
+ 177.600001n V_low
+ 177.700000n V_low
+ 177.700001n V_low
+ 177.800000n V_low
+ 177.800001n V_low
+ 177.900000n V_low
+ 177.900001n V_low
+ 178.000000n V_low
+ 178.000001n V_low
+ 178.100000n V_low
+ 178.100001n V_low
+ 178.200000n V_low
+ 178.200001n V_low
+ 178.300000n V_low
+ 178.300001n V_low
+ 178.400000n V_low
+ 178.400001n V_low
+ 178.500000n V_low
+ 178.500001n V_low
+ 178.600000n V_low
+ 178.600001n V_low
+ 178.700000n V_low
+ 178.700001n V_low
+ 178.800000n V_low
+ 178.800001n V_low
+ 178.900000n V_low
+ 178.900001n V_low
+ 179.000000n V_low
+ 179.000001n V_low
+ 179.100000n V_low
+ 179.100001n V_low
+ 179.200000n V_low
+ 179.200001n V_low
+ 179.300000n V_low
+ 179.300001n V_low
+ 179.400000n V_low
+ 179.400001n V_low
+ 179.500000n V_low
+ 179.500001n V_low
+ 179.600000n V_low
+ 179.600001n V_low
+ 179.700000n V_low
+ 179.700001n V_low
+ 179.800000n V_low
+ 179.800001n V_low
+ 179.900000n V_low
+ 179.900001n V_low
+ 180.000000n V_low
+ 180.000001n V_hig
+ 180.100000n V_hig
+ 180.100001n V_hig
+ 180.200000n V_hig
+ 180.200001n V_hig
+ 180.300000n V_hig
+ 180.300001n V_hig
+ 180.400000n V_hig
+ 180.400001n V_hig
+ 180.500000n V_hig
+ 180.500001n V_hig
+ 180.600000n V_hig
+ 180.600001n V_hig
+ 180.700000n V_hig
+ 180.700001n V_hig
+ 180.800000n V_hig
+ 180.800001n V_hig
+ 180.900000n V_hig
+ 180.900001n V_hig
+ 181.000000n V_hig
+ 181.000001n V_hig
+ 181.100000n V_hig
+ 181.100001n V_hig
+ 181.200000n V_hig
+ 181.200001n V_hig
+ 181.300000n V_hig
+ 181.300001n V_hig
+ 181.400000n V_hig
+ 181.400001n V_hig
+ 181.500000n V_hig
+ 181.500001n V_hig
+ 181.600000n V_hig
+ 181.600001n V_hig
+ 181.700000n V_hig
+ 181.700001n V_hig
+ 181.800000n V_hig
+ 181.800001n V_hig
+ 181.900000n V_hig
+ 181.900001n V_hig
+ 182.000000n V_hig
+ 182.000001n V_low
+ 182.100000n V_low
+ 182.100001n V_low
+ 182.200000n V_low
+ 182.200001n V_low
+ 182.300000n V_low
+ 182.300001n V_low
+ 182.400000n V_low
+ 182.400001n V_low
+ 182.500000n V_low
+ 182.500001n V_low
+ 182.600000n V_low
+ 182.600001n V_low
+ 182.700000n V_low
+ 182.700001n V_low
+ 182.800000n V_low
+ 182.800001n V_low
+ 182.900000n V_low
+ 182.900001n V_low
+ 183.000000n V_low
+ 183.000001n V_hig
+ 183.100000n V_hig
+ 183.100001n V_hig
+ 183.200000n V_hig
+ 183.200001n V_hig
+ 183.300000n V_hig
+ 183.300001n V_hig
+ 183.400000n V_hig
+ 183.400001n V_hig
+ 183.500000n V_hig
+ 183.500001n V_hig
+ 183.600000n V_hig
+ 183.600001n V_hig
+ 183.700000n V_hig
+ 183.700001n V_hig
+ 183.800000n V_hig
+ 183.800001n V_hig
+ 183.900000n V_hig
+ 183.900001n V_hig
+ 184.000000n V_hig
+ 184.000001n V_hig
+ 184.100000n V_hig
+ 184.100001n V_hig
+ 184.200000n V_hig
+ 184.200001n V_hig
+ 184.300000n V_hig
+ 184.300001n V_hig
+ 184.400000n V_hig
+ 184.400001n V_hig
+ 184.500000n V_hig
+ 184.500001n V_hig
+ 184.600000n V_hig
+ 184.600001n V_hig
+ 184.700000n V_hig
+ 184.700001n V_hig
+ 184.800000n V_hig
+ 184.800001n V_hig
+ 184.900000n V_hig
+ 184.900001n V_hig
+ 185.000000n V_hig
+ 185.000001n V_hig
+ 185.100000n V_hig
+ 185.100001n V_hig
+ 185.200000n V_hig
+ 185.200001n V_hig
+ 185.300000n V_hig
+ 185.300001n V_hig
+ 185.400000n V_hig
+ 185.400001n V_hig
+ 185.500000n V_hig
+ 185.500001n V_hig
+ 185.600000n V_hig
+ 185.600001n V_hig
+ 185.700000n V_hig
+ 185.700001n V_hig
+ 185.800000n V_hig
+ 185.800001n V_hig
+ 185.900000n V_hig
+ 185.900001n V_hig
+ 186.000000n V_hig
+ 186.000001n V_low
+ 186.100000n V_low
+ 186.100001n V_low
+ 186.200000n V_low
+ 186.200001n V_low
+ 186.300000n V_low
+ 186.300001n V_low
+ 186.400000n V_low
+ 186.400001n V_low
+ 186.500000n V_low
+ 186.500001n V_low
+ 186.600000n V_low
+ 186.600001n V_low
+ 186.700000n V_low
+ 186.700001n V_low
+ 186.800000n V_low
+ 186.800001n V_low
+ 186.900000n V_low
+ 186.900001n V_low
+ 187.000000n V_low
+ 187.000001n V_hig
+ 187.100000n V_hig
+ 187.100001n V_hig
+ 187.200000n V_hig
+ 187.200001n V_hig
+ 187.300000n V_hig
+ 187.300001n V_hig
+ 187.400000n V_hig
+ 187.400001n V_hig
+ 187.500000n V_hig
+ 187.500001n V_hig
+ 187.600000n V_hig
+ 187.600001n V_hig
+ 187.700000n V_hig
+ 187.700001n V_hig
+ 187.800000n V_hig
+ 187.800001n V_hig
+ 187.900000n V_hig
+ 187.900001n V_hig
+ 188.000000n V_hig
+ 188.000001n V_hig
+ 188.100000n V_hig
+ 188.100001n V_hig
+ 188.200000n V_hig
+ 188.200001n V_hig
+ 188.300000n V_hig
+ 188.300001n V_hig
+ 188.400000n V_hig
+ 188.400001n V_hig
+ 188.500000n V_hig
+ 188.500001n V_hig
+ 188.600000n V_hig
+ 188.600001n V_hig
+ 188.700000n V_hig
+ 188.700001n V_hig
+ 188.800000n V_hig
+ 188.800001n V_hig
+ 188.900000n V_hig
+ 188.900001n V_hig
+ 189.000000n V_hig
+ 189.000001n V_low
+ 189.100000n V_low
+ 189.100001n V_low
+ 189.200000n V_low
+ 189.200001n V_low
+ 189.300000n V_low
+ 189.300001n V_low
+ 189.400000n V_low
+ 189.400001n V_low
+ 189.500000n V_low
+ 189.500001n V_low
+ 189.600000n V_low
+ 189.600001n V_low
+ 189.700000n V_low
+ 189.700001n V_low
+ 189.800000n V_low
+ 189.800001n V_low
+ 189.900000n V_low
+ 189.900001n V_low
+ 190.000000n V_low
+ 190.000001n V_hig
+ 190.100000n V_hig
+ 190.100001n V_hig
+ 190.200000n V_hig
+ 190.200001n V_hig
+ 190.300000n V_hig
+ 190.300001n V_hig
+ 190.400000n V_hig
+ 190.400001n V_hig
+ 190.500000n V_hig
+ 190.500001n V_hig
+ 190.600000n V_hig
+ 190.600001n V_hig
+ 190.700000n V_hig
+ 190.700001n V_hig
+ 190.800000n V_hig
+ 190.800001n V_hig
+ 190.900000n V_hig
+ 190.900001n V_hig
+ 191.000000n V_hig
+ 191.000001n V_hig
+ 191.100000n V_hig
+ 191.100001n V_hig
+ 191.200000n V_hig
+ 191.200001n V_hig
+ 191.300000n V_hig
+ 191.300001n V_hig
+ 191.400000n V_hig
+ 191.400001n V_hig
+ 191.500000n V_hig
+ 191.500001n V_hig
+ 191.600000n V_hig
+ 191.600001n V_hig
+ 191.700000n V_hig
+ 191.700001n V_hig
+ 191.800000n V_hig
+ 191.800001n V_hig
+ 191.900000n V_hig
+ 191.900001n V_hig
+ 192.000000n V_hig
+ 192.000001n V_hig
+ 192.100000n V_hig
+ 192.100001n V_hig
+ 192.200000n V_hig
+ 192.200001n V_hig
+ 192.300000n V_hig
+ 192.300001n V_hig
+ 192.400000n V_hig
+ 192.400001n V_hig
+ 192.500000n V_hig
+ 192.500001n V_hig
+ 192.600000n V_hig
+ 192.600001n V_hig
+ 192.700000n V_hig
+ 192.700001n V_hig
+ 192.800000n V_hig
+ 192.800001n V_hig
+ 192.900000n V_hig
+ 192.900001n V_hig
+ 193.000000n V_hig
+ 193.000001n V_hig
+ 193.100000n V_hig
+ 193.100001n V_hig
+ 193.200000n V_hig
+ 193.200001n V_hig
+ 193.300000n V_hig
+ 193.300001n V_hig
+ 193.400000n V_hig
+ 193.400001n V_hig
+ 193.500000n V_hig
+ 193.500001n V_hig
+ 193.600000n V_hig
+ 193.600001n V_hig
+ 193.700000n V_hig
+ 193.700001n V_hig
+ 193.800000n V_hig
+ 193.800001n V_hig
+ 193.900000n V_hig
+ 193.900001n V_hig
+ 194.000000n V_hig
+ 194.000001n V_low
+ 194.100000n V_low
+ 194.100001n V_low
+ 194.200000n V_low
+ 194.200001n V_low
+ 194.300000n V_low
+ 194.300001n V_low
+ 194.400000n V_low
+ 194.400001n V_low
+ 194.500000n V_low
+ 194.500001n V_low
+ 194.600000n V_low
+ 194.600001n V_low
+ 194.700000n V_low
+ 194.700001n V_low
+ 194.800000n V_low
+ 194.800001n V_low
+ 194.900000n V_low
+ 194.900001n V_low
+ 195.000000n V_low
+ 195.000001n V_hig
+ 195.100000n V_hig
+ 195.100001n V_hig
+ 195.200000n V_hig
+ 195.200001n V_hig
+ 195.300000n V_hig
+ 195.300001n V_hig
+ 195.400000n V_hig
+ 195.400001n V_hig
+ 195.500000n V_hig
+ 195.500001n V_hig
+ 195.600000n V_hig
+ 195.600001n V_hig
+ 195.700000n V_hig
+ 195.700001n V_hig
+ 195.800000n V_hig
+ 195.800001n V_hig
+ 195.900000n V_hig
+ 195.900001n V_hig
+ 196.000000n V_hig
+ 196.000001n V_hig
+ 196.100000n V_hig
+ 196.100001n V_hig
+ 196.200000n V_hig
+ 196.200001n V_hig
+ 196.300000n V_hig
+ 196.300001n V_hig
+ 196.400000n V_hig
+ 196.400001n V_hig
+ 196.500000n V_hig
+ 196.500001n V_hig
+ 196.600000n V_hig
+ 196.600001n V_hig
+ 196.700000n V_hig
+ 196.700001n V_hig
+ 196.800000n V_hig
+ 196.800001n V_hig
+ 196.900000n V_hig
+ 196.900001n V_hig
+ 197.000000n V_hig
+ 197.000001n V_hig
+ 197.100000n V_hig
+ 197.100001n V_hig
+ 197.200000n V_hig
+ 197.200001n V_hig
+ 197.300000n V_hig
+ 197.300001n V_hig
+ 197.400000n V_hig
+ 197.400001n V_hig
+ 197.500000n V_hig
+ 197.500001n V_hig
+ 197.600000n V_hig
+ 197.600001n V_hig
+ 197.700000n V_hig
+ 197.700001n V_hig
+ 197.800000n V_hig
+ 197.800001n V_hig
+ 197.900000n V_hig
+ 197.900001n V_hig
+ 198.000000n V_hig
+ 198.000001n V_hig
+ 198.100000n V_hig
+ 198.100001n V_hig
+ 198.200000n V_hig
+ 198.200001n V_hig
+ 198.300000n V_hig
+ 198.300001n V_hig
+ 198.400000n V_hig
+ 198.400001n V_hig
+ 198.500000n V_hig
+ 198.500001n V_hig
+ 198.600000n V_hig
+ 198.600001n V_hig
+ 198.700000n V_hig
+ 198.700001n V_hig
+ 198.800000n V_hig
+ 198.800001n V_hig
+ 198.900000n V_hig
+ 198.900001n V_hig
+ 199.000000n V_hig
+ 199.000001n V_low
+ 199.100000n V_low
+ 199.100001n V_low
+ 199.200000n V_low
+ 199.200001n V_low
+ 199.300000n V_low
+ 199.300001n V_low
+ 199.400000n V_low
+ 199.400001n V_low
+ 199.500000n V_low
+ 199.500001n V_low
+ 199.600000n V_low
+ 199.600001n V_low
+ 199.700000n V_low
+ 199.700001n V_low
+ 199.800000n V_low
+ 199.800001n V_low
+ 199.900000n V_low
+ 199.900001n V_low
+ 200.000000n V_low
+ 200.000001n V_low
+ 200.100000n V_low
+ 200.100001n V_low
+ 200.200000n V_low
+ 200.200001n V_low
+ 200.300000n V_low
+ 200.300001n V_low
+ 200.400000n V_low
+ 200.400001n V_low
+ 200.500000n V_low
+ 200.500001n V_low
+ 200.600000n V_low
+ 200.600001n V_low
+ 200.700000n V_low
+ 200.700001n V_low
+ 200.800000n V_low
+ 200.800001n V_low
+ 200.900000n V_low
+ 200.900001n V_low
+ 201.000000n V_low
+ 201.000001n V_low
+ 201.100000n V_low
+ 201.100001n V_low
+ 201.200000n V_low
+ 201.200001n V_low
+ 201.300000n V_low
+ 201.300001n V_low
+ 201.400000n V_low
+ 201.400001n V_low
+ 201.500000n V_low
+ 201.500001n V_low
+ 201.600000n V_low
+ 201.600001n V_low
+ 201.700000n V_low
+ 201.700001n V_low
+ 201.800000n V_low
+ 201.800001n V_low
+ 201.900000n V_low
+ 201.900001n V_low
+ 202.000000n V_low
+ 202.000001n V_hig
+ 202.100000n V_hig
+ 202.100001n V_hig
+ 202.200000n V_hig
+ 202.200001n V_hig
+ 202.300000n V_hig
+ 202.300001n V_hig
+ 202.400000n V_hig
+ 202.400001n V_hig
+ 202.500000n V_hig
+ 202.500001n V_hig
+ 202.600000n V_hig
+ 202.600001n V_hig
+ 202.700000n V_hig
+ 202.700001n V_hig
+ 202.800000n V_hig
+ 202.800001n V_hig
+ 202.900000n V_hig
+ 202.900001n V_hig
+ 203.000000n V_hig
+ 203.000001n V_low
+ 203.100000n V_low
+ 203.100001n V_low
+ 203.200000n V_low
+ 203.200001n V_low
+ 203.300000n V_low
+ 203.300001n V_low
+ 203.400000n V_low
+ 203.400001n V_low
+ 203.500000n V_low
+ 203.500001n V_low
+ 203.600000n V_low
+ 203.600001n V_low
+ 203.700000n V_low
+ 203.700001n V_low
+ 203.800000n V_low
+ 203.800001n V_low
+ 203.900000n V_low
+ 203.900001n V_low
+ 204.000000n V_low
+ 204.000001n V_hig
+ 204.100000n V_hig
+ 204.100001n V_hig
+ 204.200000n V_hig
+ 204.200001n V_hig
+ 204.300000n V_hig
+ 204.300001n V_hig
+ 204.400000n V_hig
+ 204.400001n V_hig
+ 204.500000n V_hig
+ 204.500001n V_hig
+ 204.600000n V_hig
+ 204.600001n V_hig
+ 204.700000n V_hig
+ 204.700001n V_hig
+ 204.800000n V_hig
+ 204.800001n V_hig
+ 204.900000n V_hig
+ 204.900001n V_hig
+ 205.000000n V_hig
+ 205.000001n V_low
+ 205.100000n V_low
+ 205.100001n V_low
+ 205.200000n V_low
+ 205.200001n V_low
+ 205.300000n V_low
+ 205.300001n V_low
+ 205.400000n V_low
+ 205.400001n V_low
+ 205.500000n V_low
+ 205.500001n V_low
+ 205.600000n V_low
+ 205.600001n V_low
+ 205.700000n V_low
+ 205.700001n V_low
+ 205.800000n V_low
+ 205.800001n V_low
+ 205.900000n V_low
+ 205.900001n V_low
+ 206.000000n V_low
+ 206.000001n V_hig
+ 206.100000n V_hig
+ 206.100001n V_hig
+ 206.200000n V_hig
+ 206.200001n V_hig
+ 206.300000n V_hig
+ 206.300001n V_hig
+ 206.400000n V_hig
+ 206.400001n V_hig
+ 206.500000n V_hig
+ 206.500001n V_hig
+ 206.600000n V_hig
+ 206.600001n V_hig
+ 206.700000n V_hig
+ 206.700001n V_hig
+ 206.800000n V_hig
+ 206.800001n V_hig
+ 206.900000n V_hig
+ 206.900001n V_hig
+ 207.000000n V_hig
+ 207.000001n V_low
+ 207.100000n V_low
+ 207.100001n V_low
+ 207.200000n V_low
+ 207.200001n V_low
+ 207.300000n V_low
+ 207.300001n V_low
+ 207.400000n V_low
+ 207.400001n V_low
+ 207.500000n V_low
+ 207.500001n V_low
+ 207.600000n V_low
+ 207.600001n V_low
+ 207.700000n V_low
+ 207.700001n V_low
+ 207.800000n V_low
+ 207.800001n V_low
+ 207.900000n V_low
+ 207.900001n V_low
+ 208.000000n V_low
+ 208.000001n V_hig
+ 208.100000n V_hig
+ 208.100001n V_hig
+ 208.200000n V_hig
+ 208.200001n V_hig
+ 208.300000n V_hig
+ 208.300001n V_hig
+ 208.400000n V_hig
+ 208.400001n V_hig
+ 208.500000n V_hig
+ 208.500001n V_hig
+ 208.600000n V_hig
+ 208.600001n V_hig
+ 208.700000n V_hig
+ 208.700001n V_hig
+ 208.800000n V_hig
+ 208.800001n V_hig
+ 208.900000n V_hig
+ 208.900001n V_hig
+ 209.000000n V_hig
+ 209.000001n V_low
+ 209.100000n V_low
+ 209.100001n V_low
+ 209.200000n V_low
+ 209.200001n V_low
+ 209.300000n V_low
+ 209.300001n V_low
+ 209.400000n V_low
+ 209.400001n V_low
+ 209.500000n V_low
+ 209.500001n V_low
+ 209.600000n V_low
+ 209.600001n V_low
+ 209.700000n V_low
+ 209.700001n V_low
+ 209.800000n V_low
+ 209.800001n V_low
+ 209.900000n V_low
+ 209.900001n V_low
+ 210.000000n V_low
+ 210.000001n V_hig
+ 210.100000n V_hig
+ 210.100001n V_hig
+ 210.200000n V_hig
+ 210.200001n V_hig
+ 210.300000n V_hig
+ 210.300001n V_hig
+ 210.400000n V_hig
+ 210.400001n V_hig
+ 210.500000n V_hig
+ 210.500001n V_hig
+ 210.600000n V_hig
+ 210.600001n V_hig
+ 210.700000n V_hig
+ 210.700001n V_hig
+ 210.800000n V_hig
+ 210.800001n V_hig
+ 210.900000n V_hig
+ 210.900001n V_hig
+ 211.000000n V_hig
+ 211.000001n V_low
+ 211.100000n V_low
+ 211.100001n V_low
+ 211.200000n V_low
+ 211.200001n V_low
+ 211.300000n V_low
+ 211.300001n V_low
+ 211.400000n V_low
+ 211.400001n V_low
+ 211.500000n V_low
+ 211.500001n V_low
+ 211.600000n V_low
+ 211.600001n V_low
+ 211.700000n V_low
+ 211.700001n V_low
+ 211.800000n V_low
+ 211.800001n V_low
+ 211.900000n V_low
+ 211.900001n V_low
+ 212.000000n V_low
+ 212.000001n V_low
+ 212.100000n V_low
+ 212.100001n V_low
+ 212.200000n V_low
+ 212.200001n V_low
+ 212.300000n V_low
+ 212.300001n V_low
+ 212.400000n V_low
+ 212.400001n V_low
+ 212.500000n V_low
+ 212.500001n V_low
+ 212.600000n V_low
+ 212.600001n V_low
+ 212.700000n V_low
+ 212.700001n V_low
+ 212.800000n V_low
+ 212.800001n V_low
+ 212.900000n V_low
+ 212.900001n V_low
+ 213.000000n V_low
+ 213.000001n V_low
+ 213.100000n V_low
+ 213.100001n V_low
+ 213.200000n V_low
+ 213.200001n V_low
+ 213.300000n V_low
+ 213.300001n V_low
+ 213.400000n V_low
+ 213.400001n V_low
+ 213.500000n V_low
+ 213.500001n V_low
+ 213.600000n V_low
+ 213.600001n V_low
+ 213.700000n V_low
+ 213.700001n V_low
+ 213.800000n V_low
+ 213.800001n V_low
+ 213.900000n V_low
+ 213.900001n V_low
+ 214.000000n V_low
+ 214.000001n V_hig
+ 214.100000n V_hig
+ 214.100001n V_hig
+ 214.200000n V_hig
+ 214.200001n V_hig
+ 214.300000n V_hig
+ 214.300001n V_hig
+ 214.400000n V_hig
+ 214.400001n V_hig
+ 214.500000n V_hig
+ 214.500001n V_hig
+ 214.600000n V_hig
+ 214.600001n V_hig
+ 214.700000n V_hig
+ 214.700001n V_hig
+ 214.800000n V_hig
+ 214.800001n V_hig
+ 214.900000n V_hig
+ 214.900001n V_hig
+ 215.000000n V_hig
+ 215.000001n V_hig
+ 215.100000n V_hig
+ 215.100001n V_hig
+ 215.200000n V_hig
+ 215.200001n V_hig
+ 215.300000n V_hig
+ 215.300001n V_hig
+ 215.400000n V_hig
+ 215.400001n V_hig
+ 215.500000n V_hig
+ 215.500001n V_hig
+ 215.600000n V_hig
+ 215.600001n V_hig
+ 215.700000n V_hig
+ 215.700001n V_hig
+ 215.800000n V_hig
+ 215.800001n V_hig
+ 215.900000n V_hig
+ 215.900001n V_hig
+ 216.000000n V_hig
+ 216.000001n V_low
+ 216.100000n V_low
+ 216.100001n V_low
+ 216.200000n V_low
+ 216.200001n V_low
+ 216.300000n V_low
+ 216.300001n V_low
+ 216.400000n V_low
+ 216.400001n V_low
+ 216.500000n V_low
+ 216.500001n V_low
+ 216.600000n V_low
+ 216.600001n V_low
+ 216.700000n V_low
+ 216.700001n V_low
+ 216.800000n V_low
+ 216.800001n V_low
+ 216.900000n V_low
+ 216.900001n V_low
+ 217.000000n V_low
+ 217.000001n V_hig
+ 217.100000n V_hig
+ 217.100001n V_hig
+ 217.200000n V_hig
+ 217.200001n V_hig
+ 217.300000n V_hig
+ 217.300001n V_hig
+ 217.400000n V_hig
+ 217.400001n V_hig
+ 217.500000n V_hig
+ 217.500001n V_hig
+ 217.600000n V_hig
+ 217.600001n V_hig
+ 217.700000n V_hig
+ 217.700001n V_hig
+ 217.800000n V_hig
+ 217.800001n V_hig
+ 217.900000n V_hig
+ 217.900001n V_hig
+ 218.000000n V_hig
+ 218.000001n V_low
+ 218.100000n V_low
+ 218.100001n V_low
+ 218.200000n V_low
+ 218.200001n V_low
+ 218.300000n V_low
+ 218.300001n V_low
+ 218.400000n V_low
+ 218.400001n V_low
+ 218.500000n V_low
+ 218.500001n V_low
+ 218.600000n V_low
+ 218.600001n V_low
+ 218.700000n V_low
+ 218.700001n V_low
+ 218.800000n V_low
+ 218.800001n V_low
+ 218.900000n V_low
+ 218.900001n V_low
+ 219.000000n V_low
+ 219.000001n V_hig
+ 219.100000n V_hig
+ 219.100001n V_hig
+ 219.200000n V_hig
+ 219.200001n V_hig
+ 219.300000n V_hig
+ 219.300001n V_hig
+ 219.400000n V_hig
+ 219.400001n V_hig
+ 219.500000n V_hig
+ 219.500001n V_hig
+ 219.600000n V_hig
+ 219.600001n V_hig
+ 219.700000n V_hig
+ 219.700001n V_hig
+ 219.800000n V_hig
+ 219.800001n V_hig
+ 219.900000n V_hig
+ 219.900001n V_hig
+ 220.000000n V_hig
+ 220.000001n V_low
+ 220.100000n V_low
+ 220.100001n V_low
+ 220.200000n V_low
+ 220.200001n V_low
+ 220.300000n V_low
+ 220.300001n V_low
+ 220.400000n V_low
+ 220.400001n V_low
+ 220.500000n V_low
+ 220.500001n V_low
+ 220.600000n V_low
+ 220.600001n V_low
+ 220.700000n V_low
+ 220.700001n V_low
+ 220.800000n V_low
+ 220.800001n V_low
+ 220.900000n V_low
+ 220.900001n V_low
+ 221.000000n V_low
+ 221.000001n V_low
+ 221.100000n V_low
+ 221.100001n V_low
+ 221.200000n V_low
+ 221.200001n V_low
+ 221.300000n V_low
+ 221.300001n V_low
+ 221.400000n V_low
+ 221.400001n V_low
+ 221.500000n V_low
+ 221.500001n V_low
+ 221.600000n V_low
+ 221.600001n V_low
+ 221.700000n V_low
+ 221.700001n V_low
+ 221.800000n V_low
+ 221.800001n V_low
+ 221.900000n V_low
+ 221.900001n V_low
+ 222.000000n V_low
+ 222.000001n V_low
+ 222.100000n V_low
+ 222.100001n V_low
+ 222.200000n V_low
+ 222.200001n V_low
+ 222.300000n V_low
+ 222.300001n V_low
+ 222.400000n V_low
+ 222.400001n V_low
+ 222.500000n V_low
+ 222.500001n V_low
+ 222.600000n V_low
+ 222.600001n V_low
+ 222.700000n V_low
+ 222.700001n V_low
+ 222.800000n V_low
+ 222.800001n V_low
+ 222.900000n V_low
+ 222.900001n V_low
+ 223.000000n V_low
+ 223.000001n V_low
+ 223.100000n V_low
+ 223.100001n V_low
+ 223.200000n V_low
+ 223.200001n V_low
+ 223.300000n V_low
+ 223.300001n V_low
+ 223.400000n V_low
+ 223.400001n V_low
+ 223.500000n V_low
+ 223.500001n V_low
+ 223.600000n V_low
+ 223.600001n V_low
+ 223.700000n V_low
+ 223.700001n V_low
+ 223.800000n V_low
+ 223.800001n V_low
+ 223.900000n V_low
+ 223.900001n V_low
+ 224.000000n V_low
+ 224.000001n V_hig
+ 224.100000n V_hig
+ 224.100001n V_hig
+ 224.200000n V_hig
+ 224.200001n V_hig
+ 224.300000n V_hig
+ 224.300001n V_hig
+ 224.400000n V_hig
+ 224.400001n V_hig
+ 224.500000n V_hig
+ 224.500001n V_hig
+ 224.600000n V_hig
+ 224.600001n V_hig
+ 224.700000n V_hig
+ 224.700001n V_hig
+ 224.800000n V_hig
+ 224.800001n V_hig
+ 224.900000n V_hig
+ 224.900001n V_hig
+ 225.000000n V_hig
+ 225.000001n V_low
+ 225.100000n V_low
+ 225.100001n V_low
+ 225.200000n V_low
+ 225.200001n V_low
+ 225.300000n V_low
+ 225.300001n V_low
+ 225.400000n V_low
+ 225.400001n V_low
+ 225.500000n V_low
+ 225.500001n V_low
+ 225.600000n V_low
+ 225.600001n V_low
+ 225.700000n V_low
+ 225.700001n V_low
+ 225.800000n V_low
+ 225.800001n V_low
+ 225.900000n V_low
+ 225.900001n V_low
+ 226.000000n V_low
+ 226.000001n V_low
+ 226.100000n V_low
+ 226.100001n V_low
+ 226.200000n V_low
+ 226.200001n V_low
+ 226.300000n V_low
+ 226.300001n V_low
+ 226.400000n V_low
+ 226.400001n V_low
+ 226.500000n V_low
+ 226.500001n V_low
+ 226.600000n V_low
+ 226.600001n V_low
+ 226.700000n V_low
+ 226.700001n V_low
+ 226.800000n V_low
+ 226.800001n V_low
+ 226.900000n V_low
+ 226.900001n V_low
+ 227.000000n V_low
+ 227.000001n V_hig
+ 227.100000n V_hig
+ 227.100001n V_hig
+ 227.200000n V_hig
+ 227.200001n V_hig
+ 227.300000n V_hig
+ 227.300001n V_hig
+ 227.400000n V_hig
+ 227.400001n V_hig
+ 227.500000n V_hig
+ 227.500001n V_hig
+ 227.600000n V_hig
+ 227.600001n V_hig
+ 227.700000n V_hig
+ 227.700001n V_hig
+ 227.800000n V_hig
+ 227.800001n V_hig
+ 227.900000n V_hig
+ 227.900001n V_hig
+ 228.000000n V_hig
+ 228.000001n V_low
+ 228.100000n V_low
+ 228.100001n V_low
+ 228.200000n V_low
+ 228.200001n V_low
+ 228.300000n V_low
+ 228.300001n V_low
+ 228.400000n V_low
+ 228.400001n V_low
+ 228.500000n V_low
+ 228.500001n V_low
+ 228.600000n V_low
+ 228.600001n V_low
+ 228.700000n V_low
+ 228.700001n V_low
+ 228.800000n V_low
+ 228.800001n V_low
+ 228.900000n V_low
+ 228.900001n V_low
+ 229.000000n V_low
+ 229.000001n V_low
+ 229.100000n V_low
+ 229.100001n V_low
+ 229.200000n V_low
+ 229.200001n V_low
+ 229.300000n V_low
+ 229.300001n V_low
+ 229.400000n V_low
+ 229.400001n V_low
+ 229.500000n V_low
+ 229.500001n V_low
+ 229.600000n V_low
+ 229.600001n V_low
+ 229.700000n V_low
+ 229.700001n V_low
+ 229.800000n V_low
+ 229.800001n V_low
+ 229.900000n V_low
+ 229.900001n V_low
+ 230.000000n V_low
+ 230.000001n V_low
+ 230.100000n V_low
+ 230.100001n V_low
+ 230.200000n V_low
+ 230.200001n V_low
+ 230.300000n V_low
+ 230.300001n V_low
+ 230.400000n V_low
+ 230.400001n V_low
+ 230.500000n V_low
+ 230.500001n V_low
+ 230.600000n V_low
+ 230.600001n V_low
+ 230.700000n V_low
+ 230.700001n V_low
+ 230.800000n V_low
+ 230.800001n V_low
+ 230.900000n V_low
+ 230.900001n V_low
+ 231.000000n V_low
+ 231.000001n V_hig
+ 231.100000n V_hig
+ 231.100001n V_hig
+ 231.200000n V_hig
+ 231.200001n V_hig
+ 231.300000n V_hig
+ 231.300001n V_hig
+ 231.400000n V_hig
+ 231.400001n V_hig
+ 231.500000n V_hig
+ 231.500001n V_hig
+ 231.600000n V_hig
+ 231.600001n V_hig
+ 231.700000n V_hig
+ 231.700001n V_hig
+ 231.800000n V_hig
+ 231.800001n V_hig
+ 231.900000n V_hig
+ 231.900001n V_hig
+ 232.000000n V_hig
+ 232.000001n V_hig
+ 232.100000n V_hig
+ 232.100001n V_hig
+ 232.200000n V_hig
+ 232.200001n V_hig
+ 232.300000n V_hig
+ 232.300001n V_hig
+ 232.400000n V_hig
+ 232.400001n V_hig
+ 232.500000n V_hig
+ 232.500001n V_hig
+ 232.600000n V_hig
+ 232.600001n V_hig
+ 232.700000n V_hig
+ 232.700001n V_hig
+ 232.800000n V_hig
+ 232.800001n V_hig
+ 232.900000n V_hig
+ 232.900001n V_hig
+ 233.000000n V_hig
+ 233.000001n V_low
+ 233.100000n V_low
+ 233.100001n V_low
+ 233.200000n V_low
+ 233.200001n V_low
+ 233.300000n V_low
+ 233.300001n V_low
+ 233.400000n V_low
+ 233.400001n V_low
+ 233.500000n V_low
+ 233.500001n V_low
+ 233.600000n V_low
+ 233.600001n V_low
+ 233.700000n V_low
+ 233.700001n V_low
+ 233.800000n V_low
+ 233.800001n V_low
+ 233.900000n V_low
+ 233.900001n V_low
+ 234.000000n V_low
+ 234.000001n V_hig
+ 234.100000n V_hig
+ 234.100001n V_hig
+ 234.200000n V_hig
+ 234.200001n V_hig
+ 234.300000n V_hig
+ 234.300001n V_hig
+ 234.400000n V_hig
+ 234.400001n V_hig
+ 234.500000n V_hig
+ 234.500001n V_hig
+ 234.600000n V_hig
+ 234.600001n V_hig
+ 234.700000n V_hig
+ 234.700001n V_hig
+ 234.800000n V_hig
+ 234.800001n V_hig
+ 234.900000n V_hig
+ 234.900001n V_hig
+ 235.000000n V_hig
+ 235.000001n V_hig
+ 235.100000n V_hig
+ 235.100001n V_hig
+ 235.200000n V_hig
+ 235.200001n V_hig
+ 235.300000n V_hig
+ 235.300001n V_hig
+ 235.400000n V_hig
+ 235.400001n V_hig
+ 235.500000n V_hig
+ 235.500001n V_hig
+ 235.600000n V_hig
+ 235.600001n V_hig
+ 235.700000n V_hig
+ 235.700001n V_hig
+ 235.800000n V_hig
+ 235.800001n V_hig
+ 235.900000n V_hig
+ 235.900001n V_hig
+ 236.000000n V_hig
+ 236.000001n V_hig
+ 236.100000n V_hig
+ 236.100001n V_hig
+ 236.200000n V_hig
+ 236.200001n V_hig
+ 236.300000n V_hig
+ 236.300001n V_hig
+ 236.400000n V_hig
+ 236.400001n V_hig
+ 236.500000n V_hig
+ 236.500001n V_hig
+ 236.600000n V_hig
+ 236.600001n V_hig
+ 236.700000n V_hig
+ 236.700001n V_hig
+ 236.800000n V_hig
+ 236.800001n V_hig
+ 236.900000n V_hig
+ 236.900001n V_hig
+ 237.000000n V_hig
+ 237.000001n V_hig
+ 237.100000n V_hig
+ 237.100001n V_hig
+ 237.200000n V_hig
+ 237.200001n V_hig
+ 237.300000n V_hig
+ 237.300001n V_hig
+ 237.400000n V_hig
+ 237.400001n V_hig
+ 237.500000n V_hig
+ 237.500001n V_hig
+ 237.600000n V_hig
+ 237.600001n V_hig
+ 237.700000n V_hig
+ 237.700001n V_hig
+ 237.800000n V_hig
+ 237.800001n V_hig
+ 237.900000n V_hig
+ 237.900001n V_hig
+ 238.000000n V_hig
+ 238.000001n V_low
+ 238.100000n V_low
+ 238.100001n V_low
+ 238.200000n V_low
+ 238.200001n V_low
+ 238.300000n V_low
+ 238.300001n V_low
+ 238.400000n V_low
+ 238.400001n V_low
+ 238.500000n V_low
+ 238.500001n V_low
+ 238.600000n V_low
+ 238.600001n V_low
+ 238.700000n V_low
+ 238.700001n V_low
+ 238.800000n V_low
+ 238.800001n V_low
+ 238.900000n V_low
+ 238.900001n V_low
+ 239.000000n V_low
+ 239.000001n V_hig
+ 239.100000n V_hig
+ 239.100001n V_hig
+ 239.200000n V_hig
+ 239.200001n V_hig
+ 239.300000n V_hig
+ 239.300001n V_hig
+ 239.400000n V_hig
+ 239.400001n V_hig
+ 239.500000n V_hig
+ 239.500001n V_hig
+ 239.600000n V_hig
+ 239.600001n V_hig
+ 239.700000n V_hig
+ 239.700001n V_hig
+ 239.800000n V_hig
+ 239.800001n V_hig
+ 239.900000n V_hig
+ 239.900001n V_hig
+ 240.000000n V_hig
+ 240.000001n V_low
+ 240.100000n V_low
+ 240.100001n V_low
+ 240.200000n V_low
+ 240.200001n V_low
+ 240.300000n V_low
+ 240.300001n V_low
+ 240.400000n V_low
+ 240.400001n V_low
+ 240.500000n V_low
+ 240.500001n V_low
+ 240.600000n V_low
+ 240.600001n V_low
+ 240.700000n V_low
+ 240.700001n V_low
+ 240.800000n V_low
+ 240.800001n V_low
+ 240.900000n V_low
+ 240.900001n V_low
+ 241.000000n V_low
+ 241.000001n V_low
+ 241.100000n V_low
+ 241.100001n V_low
+ 241.200000n V_low
+ 241.200001n V_low
+ 241.300000n V_low
+ 241.300001n V_low
+ 241.400000n V_low
+ 241.400001n V_low
+ 241.500000n V_low
+ 241.500001n V_low
+ 241.600000n V_low
+ 241.600001n V_low
+ 241.700000n V_low
+ 241.700001n V_low
+ 241.800000n V_low
+ 241.800001n V_low
+ 241.900000n V_low
+ 241.900001n V_low
+ 242.000000n V_low
+ 242.000001n V_low
+ 242.100000n V_low
+ 242.100001n V_low
+ 242.200000n V_low
+ 242.200001n V_low
+ 242.300000n V_low
+ 242.300001n V_low
+ 242.400000n V_low
+ 242.400001n V_low
+ 242.500000n V_low
+ 242.500001n V_low
+ 242.600000n V_low
+ 242.600001n V_low
+ 242.700000n V_low
+ 242.700001n V_low
+ 242.800000n V_low
+ 242.800001n V_low
+ 242.900000n V_low
+ 242.900001n V_low
+ 243.000000n V_low
+ 243.000001n V_hig
+ 243.100000n V_hig
+ 243.100001n V_hig
+ 243.200000n V_hig
+ 243.200001n V_hig
+ 243.300000n V_hig
+ 243.300001n V_hig
+ 243.400000n V_hig
+ 243.400001n V_hig
+ 243.500000n V_hig
+ 243.500001n V_hig
+ 243.600000n V_hig
+ 243.600001n V_hig
+ 243.700000n V_hig
+ 243.700001n V_hig
+ 243.800000n V_hig
+ 243.800001n V_hig
+ 243.900000n V_hig
+ 243.900001n V_hig
+ 244.000000n V_hig
+ 244.000001n V_low
+ 244.100000n V_low
+ 244.100001n V_low
+ 244.200000n V_low
+ 244.200001n V_low
+ 244.300000n V_low
+ 244.300001n V_low
+ 244.400000n V_low
+ 244.400001n V_low
+ 244.500000n V_low
+ 244.500001n V_low
+ 244.600000n V_low
+ 244.600001n V_low
+ 244.700000n V_low
+ 244.700001n V_low
+ 244.800000n V_low
+ 244.800001n V_low
+ 244.900000n V_low
+ 244.900001n V_low
+ 245.000000n V_low
+ 245.000001n V_hig
+ 245.100000n V_hig
+ 245.100001n V_hig
+ 245.200000n V_hig
+ 245.200001n V_hig
+ 245.300000n V_hig
+ 245.300001n V_hig
+ 245.400000n V_hig
+ 245.400001n V_hig
+ 245.500000n V_hig
+ 245.500001n V_hig
+ 245.600000n V_hig
+ 245.600001n V_hig
+ 245.700000n V_hig
+ 245.700001n V_hig
+ 245.800000n V_hig
+ 245.800001n V_hig
+ 245.900000n V_hig
+ 245.900001n V_hig
+ 246.000000n V_hig
+ 246.000001n V_low
+ 246.100000n V_low
+ 246.100001n V_low
+ 246.200000n V_low
+ 246.200001n V_low
+ 246.300000n V_low
+ 246.300001n V_low
+ 246.400000n V_low
+ 246.400001n V_low
+ 246.500000n V_low
+ 246.500001n V_low
+ 246.600000n V_low
+ 246.600001n V_low
+ 246.700000n V_low
+ 246.700001n V_low
+ 246.800000n V_low
+ 246.800001n V_low
+ 246.900000n V_low
+ 246.900001n V_low
+ 247.000000n V_low
+ 247.000001n V_hig
+ 247.100000n V_hig
+ 247.100001n V_hig
+ 247.200000n V_hig
+ 247.200001n V_hig
+ 247.300000n V_hig
+ 247.300001n V_hig
+ 247.400000n V_hig
+ 247.400001n V_hig
+ 247.500000n V_hig
+ 247.500001n V_hig
+ 247.600000n V_hig
+ 247.600001n V_hig
+ 247.700000n V_hig
+ 247.700001n V_hig
+ 247.800000n V_hig
+ 247.800001n V_hig
+ 247.900000n V_hig
+ 247.900001n V_hig
+ 248.000000n V_hig
+ 248.000001n V_low
+ 248.100000n V_low
+ 248.100001n V_low
+ 248.200000n V_low
+ 248.200001n V_low
+ 248.300000n V_low
+ 248.300001n V_low
+ 248.400000n V_low
+ 248.400001n V_low
+ 248.500000n V_low
+ 248.500001n V_low
+ 248.600000n V_low
+ 248.600001n V_low
+ 248.700000n V_low
+ 248.700001n V_low
+ 248.800000n V_low
+ 248.800001n V_low
+ 248.900000n V_low
+ 248.900001n V_low
+ 249.000000n V_low
+ 249.000001n V_low
+ 249.100000n V_low
+ 249.100001n V_low
+ 249.200000n V_low
+ 249.200001n V_low
+ 249.300000n V_low
+ 249.300001n V_low
+ 249.400000n V_low
+ 249.400001n V_low
+ 249.500000n V_low
+ 249.500001n V_low
+ 249.600000n V_low
+ 249.600001n V_low
+ 249.700000n V_low
+ 249.700001n V_low
+ 249.800000n V_low
+ 249.800001n V_low
+ 249.900000n V_low
+ 249.900001n V_low
+ 250.000000n V_low
+ 250.000001n V_low
+ 250.100000n V_low
+ 250.100001n V_low
+ 250.200000n V_low
+ 250.200001n V_low
+ 250.300000n V_low
+ 250.300001n V_low
+ 250.400000n V_low
+ 250.400001n V_low
+ 250.500000n V_low
+ 250.500001n V_low
+ 250.600000n V_low
+ 250.600001n V_low
+ 250.700000n V_low
+ 250.700001n V_low
+ 250.800000n V_low
+ 250.800001n V_low
+ 250.900000n V_low
+ 250.900001n V_low
+ 251.000000n V_low
+ 251.000001n V_low
+ 251.100000n V_low
+ 251.100001n V_low
+ 251.200000n V_low
+ 251.200001n V_low
+ 251.300000n V_low
+ 251.300001n V_low
+ 251.400000n V_low
+ 251.400001n V_low
+ 251.500000n V_low
+ 251.500001n V_low
+ 251.600000n V_low
+ 251.600001n V_low
+ 251.700000n V_low
+ 251.700001n V_low
+ 251.800000n V_low
+ 251.800001n V_low
+ 251.900000n V_low
+ 251.900001n V_low
+ 252.000000n V_low
+ 252.000001n V_low
+ 252.100000n V_low
+ 252.100001n V_low
+ 252.200000n V_low
+ 252.200001n V_low
+ 252.300000n V_low
+ 252.300001n V_low
+ 252.400000n V_low
+ 252.400001n V_low
+ 252.500000n V_low
+ 252.500001n V_low
+ 252.600000n V_low
+ 252.600001n V_low
+ 252.700000n V_low
+ 252.700001n V_low
+ 252.800000n V_low
+ 252.800001n V_low
+ 252.900000n V_low
+ 252.900001n V_low
+ 253.000000n V_low
+ 253.000001n V_hig
+ 253.100000n V_hig
+ 253.100001n V_hig
+ 253.200000n V_hig
+ 253.200001n V_hig
+ 253.300000n V_hig
+ 253.300001n V_hig
+ 253.400000n V_hig
+ 253.400001n V_hig
+ 253.500000n V_hig
+ 253.500001n V_hig
+ 253.600000n V_hig
+ 253.600001n V_hig
+ 253.700000n V_hig
+ 253.700001n V_hig
+ 253.800000n V_hig
+ 253.800001n V_hig
+ 253.900000n V_hig
+ 253.900001n V_hig
+ 254.000000n V_hig
+ 254.000001n V_low
+ 254.100000n V_low
+ 254.100001n V_low
+ 254.200000n V_low
+ 254.200001n V_low
+ 254.300000n V_low
+ 254.300001n V_low
+ 254.400000n V_low
+ 254.400001n V_low
+ 254.500000n V_low
+ 254.500001n V_low
+ 254.600000n V_low
+ 254.600001n V_low
+ 254.700000n V_low
+ 254.700001n V_low
+ 254.800000n V_low
+ 254.800001n V_low
+ 254.900000n V_low
+ 254.900001n V_low
+ 255.000000n V_low
+ 255.000001n V_low
+ 255.100000n V_low
+ 255.100001n V_low
+ 255.200000n V_low
+ 255.200001n V_low
+ 255.300000n V_low
+ 255.300001n V_low
+ 255.400000n V_low
+ 255.400001n V_low
+ 255.500000n V_low
+ 255.500001n V_low
+ 255.600000n V_low
+ 255.600001n V_low
+ 255.700000n V_low
+ 255.700001n V_low
+ 255.800000n V_low
+ 255.800001n V_low
+ 255.900000n V_low
+ 255.900001n V_low
+ 256.000000n V_low
+ 256.000001n V_hig
+ 256.100000n V_hig
+ 256.100001n V_hig
+ 256.200000n V_hig
+ 256.200001n V_hig
+ 256.300000n V_hig
+ 256.300001n V_hig
+ 256.400000n V_hig
+ 256.400001n V_hig
+ 256.500000n V_hig
+ 256.500001n V_hig
+ 256.600000n V_hig
+ 256.600001n V_hig
+ 256.700000n V_hig
+ 256.700001n V_hig
+ 256.800000n V_hig
+ 256.800001n V_hig
+ 256.900000n V_hig
+ 256.900001n V_hig
+ 257.000000n V_hig
+ 257.000001n V_low
+ 257.100000n V_low
+ 257.100001n V_low
+ 257.200000n V_low
+ 257.200001n V_low
+ 257.300000n V_low
+ 257.300001n V_low
+ 257.400000n V_low
+ 257.400001n V_low
+ 257.500000n V_low
+ 257.500001n V_low
+ 257.600000n V_low
+ 257.600001n V_low
+ 257.700000n V_low
+ 257.700001n V_low
+ 257.800000n V_low
+ 257.800001n V_low
+ 257.900000n V_low
+ 257.900001n V_low
+ 258.000000n V_low
+ 258.000001n V_low
+ 258.100000n V_low
+ 258.100001n V_low
+ 258.200000n V_low
+ 258.200001n V_low
+ 258.300000n V_low
+ 258.300001n V_low
+ 258.400000n V_low
+ 258.400001n V_low
+ 258.500000n V_low
+ 258.500001n V_low
+ 258.600000n V_low
+ 258.600001n V_low
+ 258.700000n V_low
+ 258.700001n V_low
+ 258.800000n V_low
+ 258.800001n V_low
+ 258.900000n V_low
+ 258.900001n V_low
+ 259.000000n V_low
+ 259.000001n V_hig
+ 259.100000n V_hig
+ 259.100001n V_hig
+ 259.200000n V_hig
+ 259.200001n V_hig
+ 259.300000n V_hig
+ 259.300001n V_hig
+ 259.400000n V_hig
+ 259.400001n V_hig
+ 259.500000n V_hig
+ 259.500001n V_hig
+ 259.600000n V_hig
+ 259.600001n V_hig
+ 259.700000n V_hig
+ 259.700001n V_hig
+ 259.800000n V_hig
+ 259.800001n V_hig
+ 259.900000n V_hig
+ 259.900001n V_hig
+ 260.000000n V_hig
+ 260.000001n V_low
+ 260.100000n V_low
+ 260.100001n V_low
+ 260.200000n V_low
+ 260.200001n V_low
+ 260.300000n V_low
+ 260.300001n V_low
+ 260.400000n V_low
+ 260.400001n V_low
+ 260.500000n V_low
+ 260.500001n V_low
+ 260.600000n V_low
+ 260.600001n V_low
+ 260.700000n V_low
+ 260.700001n V_low
+ 260.800000n V_low
+ 260.800001n V_low
+ 260.900000n V_low
+ 260.900001n V_low
+ 261.000000n V_low
+ 261.000001n V_low
+ 261.100000n V_low
+ 261.100001n V_low
+ 261.200000n V_low
+ 261.200001n V_low
+ 261.300000n V_low
+ 261.300001n V_low
+ 261.400000n V_low
+ 261.400001n V_low
+ 261.500000n V_low
+ 261.500001n V_low
+ 261.600000n V_low
+ 261.600001n V_low
+ 261.700000n V_low
+ 261.700001n V_low
+ 261.800000n V_low
+ 261.800001n V_low
+ 261.900000n V_low
+ 261.900001n V_low
+ 262.000000n V_low
+ 262.000001n V_hig
+ 262.100000n V_hig
+ 262.100001n V_hig
+ 262.200000n V_hig
+ 262.200001n V_hig
+ 262.300000n V_hig
+ 262.300001n V_hig
+ 262.400000n V_hig
+ 262.400001n V_hig
+ 262.500000n V_hig
+ 262.500001n V_hig
+ 262.600000n V_hig
+ 262.600001n V_hig
+ 262.700000n V_hig
+ 262.700001n V_hig
+ 262.800000n V_hig
+ 262.800001n V_hig
+ 262.900000n V_hig
+ 262.900001n V_hig
+ 263.000000n V_hig
+ 263.000001n V_hig
+ 263.100000n V_hig
+ 263.100001n V_hig
+ 263.200000n V_hig
+ 263.200001n V_hig
+ 263.300000n V_hig
+ 263.300001n V_hig
+ 263.400000n V_hig
+ 263.400001n V_hig
+ 263.500000n V_hig
+ 263.500001n V_hig
+ 263.600000n V_hig
+ 263.600001n V_hig
+ 263.700000n V_hig
+ 263.700001n V_hig
+ 263.800000n V_hig
+ 263.800001n V_hig
+ 263.900000n V_hig
+ 263.900001n V_hig
+ 264.000000n V_hig
+ 264.000001n V_hig
+ 264.100000n V_hig
+ 264.100001n V_hig
+ 264.200000n V_hig
+ 264.200001n V_hig
+ 264.300000n V_hig
+ 264.300001n V_hig
+ 264.400000n V_hig
+ 264.400001n V_hig
+ 264.500000n V_hig
+ 264.500001n V_hig
+ 264.600000n V_hig
+ 264.600001n V_hig
+ 264.700000n V_hig
+ 264.700001n V_hig
+ 264.800000n V_hig
+ 264.800001n V_hig
+ 264.900000n V_hig
+ 264.900001n V_hig
+ 265.000000n V_hig
+ 265.000001n V_low
+ 265.100000n V_low
+ 265.100001n V_low
+ 265.200000n V_low
+ 265.200001n V_low
+ 265.300000n V_low
+ 265.300001n V_low
+ 265.400000n V_low
+ 265.400001n V_low
+ 265.500000n V_low
+ 265.500001n V_low
+ 265.600000n V_low
+ 265.600001n V_low
+ 265.700000n V_low
+ 265.700001n V_low
+ 265.800000n V_low
+ 265.800001n V_low
+ 265.900000n V_low
+ 265.900001n V_low
+ 266.000000n V_low
+ 266.000001n V_hig
+ 266.100000n V_hig
+ 266.100001n V_hig
+ 266.200000n V_hig
+ 266.200001n V_hig
+ 266.300000n V_hig
+ 266.300001n V_hig
+ 266.400000n V_hig
+ 266.400001n V_hig
+ 266.500000n V_hig
+ 266.500001n V_hig
+ 266.600000n V_hig
+ 266.600001n V_hig
+ 266.700000n V_hig
+ 266.700001n V_hig
+ 266.800000n V_hig
+ 266.800001n V_hig
+ 266.900000n V_hig
+ 266.900001n V_hig
+ 267.000000n V_hig
+ 267.000001n V_hig
+ 267.100000n V_hig
+ 267.100001n V_hig
+ 267.200000n V_hig
+ 267.200001n V_hig
+ 267.300000n V_hig
+ 267.300001n V_hig
+ 267.400000n V_hig
+ 267.400001n V_hig
+ 267.500000n V_hig
+ 267.500001n V_hig
+ 267.600000n V_hig
+ 267.600001n V_hig
+ 267.700000n V_hig
+ 267.700001n V_hig
+ 267.800000n V_hig
+ 267.800001n V_hig
+ 267.900000n V_hig
+ 267.900001n V_hig
+ 268.000000n V_hig
+ 268.000001n V_hig
+ 268.100000n V_hig
+ 268.100001n V_hig
+ 268.200000n V_hig
+ 268.200001n V_hig
+ 268.300000n V_hig
+ 268.300001n V_hig
+ 268.400000n V_hig
+ 268.400001n V_hig
+ 268.500000n V_hig
+ 268.500001n V_hig
+ 268.600000n V_hig
+ 268.600001n V_hig
+ 268.700000n V_hig
+ 268.700001n V_hig
+ 268.800000n V_hig
+ 268.800001n V_hig
+ 268.900000n V_hig
+ 268.900001n V_hig
+ 269.000000n V_hig
+ 269.000001n V_hig
+ 269.100000n V_hig
+ 269.100001n V_hig
+ 269.200000n V_hig
+ 269.200001n V_hig
+ 269.300000n V_hig
+ 269.300001n V_hig
+ 269.400000n V_hig
+ 269.400001n V_hig
+ 269.500000n V_hig
+ 269.500001n V_hig
+ 269.600000n V_hig
+ 269.600001n V_hig
+ 269.700000n V_hig
+ 269.700001n V_hig
+ 269.800000n V_hig
+ 269.800001n V_hig
+ 269.900000n V_hig
+ 269.900001n V_hig
+ 270.000000n V_hig
+ 270.000001n V_low
+ 270.100000n V_low
+ 270.100001n V_low
+ 270.200000n V_low
+ 270.200001n V_low
+ 270.300000n V_low
+ 270.300001n V_low
+ 270.400000n V_low
+ 270.400001n V_low
+ 270.500000n V_low
+ 270.500001n V_low
+ 270.600000n V_low
+ 270.600001n V_low
+ 270.700000n V_low
+ 270.700001n V_low
+ 270.800000n V_low
+ 270.800001n V_low
+ 270.900000n V_low
+ 270.900001n V_low
+ 271.000000n V_low
+ 271.000001n V_hig
+ 271.100000n V_hig
+ 271.100001n V_hig
+ 271.200000n V_hig
+ 271.200001n V_hig
+ 271.300000n V_hig
+ 271.300001n V_hig
+ 271.400000n V_hig
+ 271.400001n V_hig
+ 271.500000n V_hig
+ 271.500001n V_hig
+ 271.600000n V_hig
+ 271.600001n V_hig
+ 271.700000n V_hig
+ 271.700001n V_hig
+ 271.800000n V_hig
+ 271.800001n V_hig
+ 271.900000n V_hig
+ 271.900001n V_hig
+ 272.000000n V_hig
+ 272.000001n V_low
+ 272.100000n V_low
+ 272.100001n V_low
+ 272.200000n V_low
+ 272.200001n V_low
+ 272.300000n V_low
+ 272.300001n V_low
+ 272.400000n V_low
+ 272.400001n V_low
+ 272.500000n V_low
+ 272.500001n V_low
+ 272.600000n V_low
+ 272.600001n V_low
+ 272.700000n V_low
+ 272.700001n V_low
+ 272.800000n V_low
+ 272.800001n V_low
+ 272.900000n V_low
+ 272.900001n V_low
+ 273.000000n V_low
+ 273.000001n V_low
+ 273.100000n V_low
+ 273.100001n V_low
+ 273.200000n V_low
+ 273.200001n V_low
+ 273.300000n V_low
+ 273.300001n V_low
+ 273.400000n V_low
+ 273.400001n V_low
+ 273.500000n V_low
+ 273.500001n V_low
+ 273.600000n V_low
+ 273.600001n V_low
+ 273.700000n V_low
+ 273.700001n V_low
+ 273.800000n V_low
+ 273.800001n V_low
+ 273.900000n V_low
+ 273.900001n V_low
+ 274.000000n V_low
+ 274.000001n V_hig
+ 274.100000n V_hig
+ 274.100001n V_hig
+ 274.200000n V_hig
+ 274.200001n V_hig
+ 274.300000n V_hig
+ 274.300001n V_hig
+ 274.400000n V_hig
+ 274.400001n V_hig
+ 274.500000n V_hig
+ 274.500001n V_hig
+ 274.600000n V_hig
+ 274.600001n V_hig
+ 274.700000n V_hig
+ 274.700001n V_hig
+ 274.800000n V_hig
+ 274.800001n V_hig
+ 274.900000n V_hig
+ 274.900001n V_hig
+ 275.000000n V_hig
+ 275.000001n V_low
+ 275.100000n V_low
+ 275.100001n V_low
+ 275.200000n V_low
+ 275.200001n V_low
+ 275.300000n V_low
+ 275.300001n V_low
+ 275.400000n V_low
+ 275.400001n V_low
+ 275.500000n V_low
+ 275.500001n V_low
+ 275.600000n V_low
+ 275.600001n V_low
+ 275.700000n V_low
+ 275.700001n V_low
+ 275.800000n V_low
+ 275.800001n V_low
+ 275.900000n V_low
+ 275.900001n V_low
+ 276.000000n V_low
+ 276.000001n V_hig
+ 276.100000n V_hig
+ 276.100001n V_hig
+ 276.200000n V_hig
+ 276.200001n V_hig
+ 276.300000n V_hig
+ 276.300001n V_hig
+ 276.400000n V_hig
+ 276.400001n V_hig
+ 276.500000n V_hig
+ 276.500001n V_hig
+ 276.600000n V_hig
+ 276.600001n V_hig
+ 276.700000n V_hig
+ 276.700001n V_hig
+ 276.800000n V_hig
+ 276.800001n V_hig
+ 276.900000n V_hig
+ 276.900001n V_hig
+ 277.000000n V_hig
+ 277.000001n V_low
+ 277.100000n V_low
+ 277.100001n V_low
+ 277.200000n V_low
+ 277.200001n V_low
+ 277.300000n V_low
+ 277.300001n V_low
+ 277.400000n V_low
+ 277.400001n V_low
+ 277.500000n V_low
+ 277.500001n V_low
+ 277.600000n V_low
+ 277.600001n V_low
+ 277.700000n V_low
+ 277.700001n V_low
+ 277.800000n V_low
+ 277.800001n V_low
+ 277.900000n V_low
+ 277.900001n V_low
+ 278.000000n V_low
+ 278.000001n V_low
+ 278.100000n V_low
+ 278.100001n V_low
+ 278.200000n V_low
+ 278.200001n V_low
+ 278.300000n V_low
+ 278.300001n V_low
+ 278.400000n V_low
+ 278.400001n V_low
+ 278.500000n V_low
+ 278.500001n V_low
+ 278.600000n V_low
+ 278.600001n V_low
+ 278.700000n V_low
+ 278.700001n V_low
+ 278.800000n V_low
+ 278.800001n V_low
+ 278.900000n V_low
+ 278.900001n V_low
+ 279.000000n V_low
+ 279.000001n V_low
+ 279.100000n V_low
+ 279.100001n V_low
+ 279.200000n V_low
+ 279.200001n V_low
+ 279.300000n V_low
+ 279.300001n V_low
+ 279.400000n V_low
+ 279.400001n V_low
+ 279.500000n V_low
+ 279.500001n V_low
+ 279.600000n V_low
+ 279.600001n V_low
+ 279.700000n V_low
+ 279.700001n V_low
+ 279.800000n V_low
+ 279.800001n V_low
+ 279.900000n V_low
+ 279.900001n V_low
+ 280.000000n V_low
+ 280.000001n V_hig
+ 280.100000n V_hig
+ 280.100001n V_hig
+ 280.200000n V_hig
+ 280.200001n V_hig
+ 280.300000n V_hig
+ 280.300001n V_hig
+ 280.400000n V_hig
+ 280.400001n V_hig
+ 280.500000n V_hig
+ 280.500001n V_hig
+ 280.600000n V_hig
+ 280.600001n V_hig
+ 280.700000n V_hig
+ 280.700001n V_hig
+ 280.800000n V_hig
+ 280.800001n V_hig
+ 280.900000n V_hig
+ 280.900001n V_hig
+ 281.000000n V_hig
+ 281.000001n V_hig
+ 281.100000n V_hig
+ 281.100001n V_hig
+ 281.200000n V_hig
+ 281.200001n V_hig
+ 281.300000n V_hig
+ 281.300001n V_hig
+ 281.400000n V_hig
+ 281.400001n V_hig
+ 281.500000n V_hig
+ 281.500001n V_hig
+ 281.600000n V_hig
+ 281.600001n V_hig
+ 281.700000n V_hig
+ 281.700001n V_hig
+ 281.800000n V_hig
+ 281.800001n V_hig
+ 281.900000n V_hig
+ 281.900001n V_hig
+ 282.000000n V_hig
+ 282.000001n V_hig
+ 282.100000n V_hig
+ 282.100001n V_hig
+ 282.200000n V_hig
+ 282.200001n V_hig
+ 282.300000n V_hig
+ 282.300001n V_hig
+ 282.400000n V_hig
+ 282.400001n V_hig
+ 282.500000n V_hig
+ 282.500001n V_hig
+ 282.600000n V_hig
+ 282.600001n V_hig
+ 282.700000n V_hig
+ 282.700001n V_hig
+ 282.800000n V_hig
+ 282.800001n V_hig
+ 282.900000n V_hig
+ 282.900001n V_hig
+ 283.000000n V_hig
+ 283.000001n V_hig
+ 283.100000n V_hig
+ 283.100001n V_hig
+ 283.200000n V_hig
+ 283.200001n V_hig
+ 283.300000n V_hig
+ 283.300001n V_hig
+ 283.400000n V_hig
+ 283.400001n V_hig
+ 283.500000n V_hig
+ 283.500001n V_hig
+ 283.600000n V_hig
+ 283.600001n V_hig
+ 283.700000n V_hig
+ 283.700001n V_hig
+ 283.800000n V_hig
+ 283.800001n V_hig
+ 283.900000n V_hig
+ 283.900001n V_hig
+ 284.000000n V_hig
+ 284.000001n V_hig
+ 284.100000n V_hig
+ 284.100001n V_hig
+ 284.200000n V_hig
+ 284.200001n V_hig
+ 284.300000n V_hig
+ 284.300001n V_hig
+ 284.400000n V_hig
+ 284.400001n V_hig
+ 284.500000n V_hig
+ 284.500001n V_hig
+ 284.600000n V_hig
+ 284.600001n V_hig
+ 284.700000n V_hig
+ 284.700001n V_hig
+ 284.800000n V_hig
+ 284.800001n V_hig
+ 284.900000n V_hig
+ 284.900001n V_hig
+ 285.000000n V_hig
+ 285.000001n V_hig
+ 285.100000n V_hig
+ 285.100001n V_hig
+ 285.200000n V_hig
+ 285.200001n V_hig
+ 285.300000n V_hig
+ 285.300001n V_hig
+ 285.400000n V_hig
+ 285.400001n V_hig
+ 285.500000n V_hig
+ 285.500001n V_hig
+ 285.600000n V_hig
+ 285.600001n V_hig
+ 285.700000n V_hig
+ 285.700001n V_hig
+ 285.800000n V_hig
+ 285.800001n V_hig
+ 285.900000n V_hig
+ 285.900001n V_hig
+ 286.000000n V_hig
+ 286.000001n V_hig
+ 286.100000n V_hig
+ 286.100001n V_hig
+ 286.200000n V_hig
+ 286.200001n V_hig
+ 286.300000n V_hig
+ 286.300001n V_hig
+ 286.400000n V_hig
+ 286.400001n V_hig
+ 286.500000n V_hig
+ 286.500001n V_hig
+ 286.600000n V_hig
+ 286.600001n V_hig
+ 286.700000n V_hig
+ 286.700001n V_hig
+ 286.800000n V_hig
+ 286.800001n V_hig
+ 286.900000n V_hig
+ 286.900001n V_hig
+ 287.000000n V_hig
+ 287.000001n V_low
+ 287.100000n V_low
+ 287.100001n V_low
+ 287.200000n V_low
+ 287.200001n V_low
+ 287.300000n V_low
+ 287.300001n V_low
+ 287.400000n V_low
+ 287.400001n V_low
+ 287.500000n V_low
+ 287.500001n V_low
+ 287.600000n V_low
+ 287.600001n V_low
+ 287.700000n V_low
+ 287.700001n V_low
+ 287.800000n V_low
+ 287.800001n V_low
+ 287.900000n V_low
+ 287.900001n V_low
+ 288.000000n V_low
+ 288.000001n V_low
+ 288.100000n V_low
+ 288.100001n V_low
+ 288.200000n V_low
+ 288.200001n V_low
+ 288.300000n V_low
+ 288.300001n V_low
+ 288.400000n V_low
+ 288.400001n V_low
+ 288.500000n V_low
+ 288.500001n V_low
+ 288.600000n V_low
+ 288.600001n V_low
+ 288.700000n V_low
+ 288.700001n V_low
+ 288.800000n V_low
+ 288.800001n V_low
+ 288.900000n V_low
+ 288.900001n V_low
+ 289.000000n V_low
+ 289.000001n V_low
+ 289.100000n V_low
+ 289.100001n V_low
+ 289.200000n V_low
+ 289.200001n V_low
+ 289.300000n V_low
+ 289.300001n V_low
+ 289.400000n V_low
+ 289.400001n V_low
+ 289.500000n V_low
+ 289.500001n V_low
+ 289.600000n V_low
+ 289.600001n V_low
+ 289.700000n V_low
+ 289.700001n V_low
+ 289.800000n V_low
+ 289.800001n V_low
+ 289.900000n V_low
+ 289.900001n V_low
+ 290.000000n V_low
+ 290.000001n V_hig
+ 290.100000n V_hig
+ 290.100001n V_hig
+ 290.200000n V_hig
+ 290.200001n V_hig
+ 290.300000n V_hig
+ 290.300001n V_hig
+ 290.400000n V_hig
+ 290.400001n V_hig
+ 290.500000n V_hig
+ 290.500001n V_hig
+ 290.600000n V_hig
+ 290.600001n V_hig
+ 290.700000n V_hig
+ 290.700001n V_hig
+ 290.800000n V_hig
+ 290.800001n V_hig
+ 290.900000n V_hig
+ 290.900001n V_hig
+ 291.000000n V_hig
+ 291.000001n V_low
+ 291.100000n V_low
+ 291.100001n V_low
+ 291.200000n V_low
+ 291.200001n V_low
+ 291.300000n V_low
+ 291.300001n V_low
+ 291.400000n V_low
+ 291.400001n V_low
+ 291.500000n V_low
+ 291.500001n V_low
+ 291.600000n V_low
+ 291.600001n V_low
+ 291.700000n V_low
+ 291.700001n V_low
+ 291.800000n V_low
+ 291.800001n V_low
+ 291.900000n V_low
+ 291.900001n V_low
+ 292.000000n V_low
+ 292.000001n V_hig
+ 292.100000n V_hig
+ 292.100001n V_hig
+ 292.200000n V_hig
+ 292.200001n V_hig
+ 292.300000n V_hig
+ 292.300001n V_hig
+ 292.400000n V_hig
+ 292.400001n V_hig
+ 292.500000n V_hig
+ 292.500001n V_hig
+ 292.600000n V_hig
+ 292.600001n V_hig
+ 292.700000n V_hig
+ 292.700001n V_hig
+ 292.800000n V_hig
+ 292.800001n V_hig
+ 292.900000n V_hig
+ 292.900001n V_hig
+ 293.000000n V_hig
+ 293.000001n V_hig
+ 293.100000n V_hig
+ 293.100001n V_hig
+ 293.200000n V_hig
+ 293.200001n V_hig
+ 293.300000n V_hig
+ 293.300001n V_hig
+ 293.400000n V_hig
+ 293.400001n V_hig
+ 293.500000n V_hig
+ 293.500001n V_hig
+ 293.600000n V_hig
+ 293.600001n V_hig
+ 293.700000n V_hig
+ 293.700001n V_hig
+ 293.800000n V_hig
+ 293.800001n V_hig
+ 293.900000n V_hig
+ 293.900001n V_hig
+ 294.000000n V_hig
+ 294.000001n V_low
+ 294.100000n V_low
+ 294.100001n V_low
+ 294.200000n V_low
+ 294.200001n V_low
+ 294.300000n V_low
+ 294.300001n V_low
+ 294.400000n V_low
+ 294.400001n V_low
+ 294.500000n V_low
+ 294.500001n V_low
+ 294.600000n V_low
+ 294.600001n V_low
+ 294.700000n V_low
+ 294.700001n V_low
+ 294.800000n V_low
+ 294.800001n V_low
+ 294.900000n V_low
+ 294.900001n V_low
+ 295.000000n V_low
+ 295.000001n V_low
+ 295.100000n V_low
+ 295.100001n V_low
+ 295.200000n V_low
+ 295.200001n V_low
+ 295.300000n V_low
+ 295.300001n V_low
+ 295.400000n V_low
+ 295.400001n V_low
+ 295.500000n V_low
+ 295.500001n V_low
+ 295.600000n V_low
+ 295.600001n V_low
+ 295.700000n V_low
+ 295.700001n V_low
+ 295.800000n V_low
+ 295.800001n V_low
+ 295.900000n V_low
+ 295.900001n V_low
+ 296.000000n V_low
+ 296.000001n V_hig
+ 296.100000n V_hig
+ 296.100001n V_hig
+ 296.200000n V_hig
+ 296.200001n V_hig
+ 296.300000n V_hig
+ 296.300001n V_hig
+ 296.400000n V_hig
+ 296.400001n V_hig
+ 296.500000n V_hig
+ 296.500001n V_hig
+ 296.600000n V_hig
+ 296.600001n V_hig
+ 296.700000n V_hig
+ 296.700001n V_hig
+ 296.800000n V_hig
+ 296.800001n V_hig
+ 296.900000n V_hig
+ 296.900001n V_hig
+ 297.000000n V_hig
+ 297.000001n V_low
+ 297.100000n V_low
+ 297.100001n V_low
+ 297.200000n V_low
+ 297.200001n V_low
+ 297.300000n V_low
+ 297.300001n V_low
+ 297.400000n V_low
+ 297.400001n V_low
+ 297.500000n V_low
+ 297.500001n V_low
+ 297.600000n V_low
+ 297.600001n V_low
+ 297.700000n V_low
+ 297.700001n V_low
+ 297.800000n V_low
+ 297.800001n V_low
+ 297.900000n V_low
+ 297.900001n V_low
+ 298.000000n V_low
+ 298.000001n V_low
+ 298.100000n V_low
+ 298.100001n V_low
+ 298.200000n V_low
+ 298.200001n V_low
+ 298.300000n V_low
+ 298.300001n V_low
+ 298.400000n V_low
+ 298.400001n V_low
+ 298.500000n V_low
+ 298.500001n V_low
+ 298.600000n V_low
+ 298.600001n V_low
+ 298.700000n V_low
+ 298.700001n V_low
+ 298.800000n V_low
+ 298.800001n V_low
+ 298.900000n V_low
+ 298.900001n V_low
+ 299.000000n V_low
+ 299.000001n V_low
+ 299.100000n V_low
+ 299.100001n V_low
+ 299.200000n V_low
+ 299.200001n V_low
+ 299.300000n V_low
+ 299.300001n V_low
+ 299.400000n V_low
+ 299.400001n V_low
+ 299.500000n V_low
+ 299.500001n V_low
+ 299.600000n V_low
+ 299.600001n V_low
+ 299.700000n V_low
+ 299.700001n V_low
+ 299.800000n V_low
+ 299.800001n V_low
+ 299.900000n V_low
+ 299.900001n V_low
+ 300.000000n V_low
+ 300.000001n V_low
+ 300.100000n V_low
+ 300.100001n V_low
+ 300.200000n V_low
+ 300.200001n V_low
+ 300.300000n V_low
+ 300.300001n V_low
+ 300.400000n V_low
+ 300.400001n V_low
+ 300.500000n V_low
+ 300.500001n V_low
+ 300.600000n V_low
+ 300.600001n V_low
+ 300.700000n V_low
+ 300.700001n V_low
+ 300.800000n V_low
+ 300.800001n V_low
+ 300.900000n V_low
+ 300.900001n V_low
+ 301.000000n V_low
+ 301.000001n V_hig
+ 301.100000n V_hig
+ 301.100001n V_hig
+ 301.200000n V_hig
+ 301.200001n V_hig
+ 301.300000n V_hig
+ 301.300001n V_hig
+ 301.400000n V_hig
+ 301.400001n V_hig
+ 301.500000n V_hig
+ 301.500001n V_hig
+ 301.600000n V_hig
+ 301.600001n V_hig
+ 301.700000n V_hig
+ 301.700001n V_hig
+ 301.800000n V_hig
+ 301.800001n V_hig
+ 301.900000n V_hig
+ 301.900001n V_hig
+ 302.000000n V_hig
+ 302.000001n V_hig
+ 302.100000n V_hig
+ 302.100001n V_hig
+ 302.200000n V_hig
+ 302.200001n V_hig
+ 302.300000n V_hig
+ 302.300001n V_hig
+ 302.400000n V_hig
+ 302.400001n V_hig
+ 302.500000n V_hig
+ 302.500001n V_hig
+ 302.600000n V_hig
+ 302.600001n V_hig
+ 302.700000n V_hig
+ 302.700001n V_hig
+ 302.800000n V_hig
+ 302.800001n V_hig
+ 302.900000n V_hig
+ 302.900001n V_hig
+ 303.000000n V_hig
+ 303.000001n V_hig
+ 303.100000n V_hig
+ 303.100001n V_hig
+ 303.200000n V_hig
+ 303.200001n V_hig
+ 303.300000n V_hig
+ 303.300001n V_hig
+ 303.400000n V_hig
+ 303.400001n V_hig
+ 303.500000n V_hig
+ 303.500001n V_hig
+ 303.600000n V_hig
+ 303.600001n V_hig
+ 303.700000n V_hig
+ 303.700001n V_hig
+ 303.800000n V_hig
+ 303.800001n V_hig
+ 303.900000n V_hig
+ 303.900001n V_hig
+ 304.000000n V_hig
+ 304.000001n V_low
+ 304.100000n V_low
+ 304.100001n V_low
+ 304.200000n V_low
+ 304.200001n V_low
+ 304.300000n V_low
+ 304.300001n V_low
+ 304.400000n V_low
+ 304.400001n V_low
+ 304.500000n V_low
+ 304.500001n V_low
+ 304.600000n V_low
+ 304.600001n V_low
+ 304.700000n V_low
+ 304.700001n V_low
+ 304.800000n V_low
+ 304.800001n V_low
+ 304.900000n V_low
+ 304.900001n V_low
+ 305.000000n V_low
+ 305.000001n V_low
+ 305.100000n V_low
+ 305.100001n V_low
+ 305.200000n V_low
+ 305.200001n V_low
+ 305.300000n V_low
+ 305.300001n V_low
+ 305.400000n V_low
+ 305.400001n V_low
+ 305.500000n V_low
+ 305.500001n V_low
+ 305.600000n V_low
+ 305.600001n V_low
+ 305.700000n V_low
+ 305.700001n V_low
+ 305.800000n V_low
+ 305.800001n V_low
+ 305.900000n V_low
+ 305.900001n V_low
+ 306.000000n V_low
+ 306.000001n V_low
+ 306.100000n V_low
+ 306.100001n V_low
+ 306.200000n V_low
+ 306.200001n V_low
+ 306.300000n V_low
+ 306.300001n V_low
+ 306.400000n V_low
+ 306.400001n V_low
+ 306.500000n V_low
+ 306.500001n V_low
+ 306.600000n V_low
+ 306.600001n V_low
+ 306.700000n V_low
+ 306.700001n V_low
+ 306.800000n V_low
+ 306.800001n V_low
+ 306.900000n V_low
+ 306.900001n V_low
+ 307.000000n V_low
+ 307.000001n V_low
+ 307.100000n V_low
+ 307.100001n V_low
+ 307.200000n V_low
+ 307.200001n V_low
+ 307.300000n V_low
+ 307.300001n V_low
+ 307.400000n V_low
+ 307.400001n V_low
+ 307.500000n V_low
+ 307.500001n V_low
+ 307.600000n V_low
+ 307.600001n V_low
+ 307.700000n V_low
+ 307.700001n V_low
+ 307.800000n V_low
+ 307.800001n V_low
+ 307.900000n V_low
+ 307.900001n V_low
+ 308.000000n V_low
+ 308.000001n V_hig
+ 308.100000n V_hig
+ 308.100001n V_hig
+ 308.200000n V_hig
+ 308.200001n V_hig
+ 308.300000n V_hig
+ 308.300001n V_hig
+ 308.400000n V_hig
+ 308.400001n V_hig
+ 308.500000n V_hig
+ 308.500001n V_hig
+ 308.600000n V_hig
+ 308.600001n V_hig
+ 308.700000n V_hig
+ 308.700001n V_hig
+ 308.800000n V_hig
+ 308.800001n V_hig
+ 308.900000n V_hig
+ 308.900001n V_hig
+ 309.000000n V_hig
+ 309.000001n V_low
+ 309.100000n V_low
+ 309.100001n V_low
+ 309.200000n V_low
+ 309.200001n V_low
+ 309.300000n V_low
+ 309.300001n V_low
+ 309.400000n V_low
+ 309.400001n V_low
+ 309.500000n V_low
+ 309.500001n V_low
+ 309.600000n V_low
+ 309.600001n V_low
+ 309.700000n V_low
+ 309.700001n V_low
+ 309.800000n V_low
+ 309.800001n V_low
+ 309.900000n V_low
+ 309.900001n V_low
+ 310.000000n V_low
+ 310.000001n V_hig
+ 310.100000n V_hig
+ 310.100001n V_hig
+ 310.200000n V_hig
+ 310.200001n V_hig
+ 310.300000n V_hig
+ 310.300001n V_hig
+ 310.400000n V_hig
+ 310.400001n V_hig
+ 310.500000n V_hig
+ 310.500001n V_hig
+ 310.600000n V_hig
+ 310.600001n V_hig
+ 310.700000n V_hig
+ 310.700001n V_hig
+ 310.800000n V_hig
+ 310.800001n V_hig
+ 310.900000n V_hig
+ 310.900001n V_hig
+ 311.000000n V_hig
+ 311.000001n V_hig
+ 311.100000n V_hig
+ 311.100001n V_hig
+ 311.200000n V_hig
+ 311.200001n V_hig
+ 311.300000n V_hig
+ 311.300001n V_hig
+ 311.400000n V_hig
+ 311.400001n V_hig
+ 311.500000n V_hig
+ 311.500001n V_hig
+ 311.600000n V_hig
+ 311.600001n V_hig
+ 311.700000n V_hig
+ 311.700001n V_hig
+ 311.800000n V_hig
+ 311.800001n V_hig
+ 311.900000n V_hig
+ 311.900001n V_hig
+ 312.000000n V_hig
+ 312.000001n V_low
+ 312.100000n V_low
+ 312.100001n V_low
+ 312.200000n V_low
+ 312.200001n V_low
+ 312.300000n V_low
+ 312.300001n V_low
+ 312.400000n V_low
+ 312.400001n V_low
+ 312.500000n V_low
+ 312.500001n V_low
+ 312.600000n V_low
+ 312.600001n V_low
+ 312.700000n V_low
+ 312.700001n V_low
+ 312.800000n V_low
+ 312.800001n V_low
+ 312.900000n V_low
+ 312.900001n V_low
+ 313.000000n V_low
+ 313.000001n V_low
+ 313.100000n V_low
+ 313.100001n V_low
+ 313.200000n V_low
+ 313.200001n V_low
+ 313.300000n V_low
+ 313.300001n V_low
+ 313.400000n V_low
+ 313.400001n V_low
+ 313.500000n V_low
+ 313.500001n V_low
+ 313.600000n V_low
+ 313.600001n V_low
+ 313.700000n V_low
+ 313.700001n V_low
+ 313.800000n V_low
+ 313.800001n V_low
+ 313.900000n V_low
+ 313.900001n V_low
+ 314.000000n V_low
+ 314.000001n V_hig
+ 314.100000n V_hig
+ 314.100001n V_hig
+ 314.200000n V_hig
+ 314.200001n V_hig
+ 314.300000n V_hig
+ 314.300001n V_hig
+ 314.400000n V_hig
+ 314.400001n V_hig
+ 314.500000n V_hig
+ 314.500001n V_hig
+ 314.600000n V_hig
+ 314.600001n V_hig
+ 314.700000n V_hig
+ 314.700001n V_hig
+ 314.800000n V_hig
+ 314.800001n V_hig
+ 314.900000n V_hig
+ 314.900001n V_hig
+ 315.000000n V_hig
+ 315.000001n V_hig
+ 315.100000n V_hig
+ 315.100001n V_hig
+ 315.200000n V_hig
+ 315.200001n V_hig
+ 315.300000n V_hig
+ 315.300001n V_hig
+ 315.400000n V_hig
+ 315.400001n V_hig
+ 315.500000n V_hig
+ 315.500001n V_hig
+ 315.600000n V_hig
+ 315.600001n V_hig
+ 315.700000n V_hig
+ 315.700001n V_hig
+ 315.800000n V_hig
+ 315.800001n V_hig
+ 315.900000n V_hig
+ 315.900001n V_hig
+ 316.000000n V_hig
+ 316.000001n V_low
+ 316.100000n V_low
+ 316.100001n V_low
+ 316.200000n V_low
+ 316.200001n V_low
+ 316.300000n V_low
+ 316.300001n V_low
+ 316.400000n V_low
+ 316.400001n V_low
+ 316.500000n V_low
+ 316.500001n V_low
+ 316.600000n V_low
+ 316.600001n V_low
+ 316.700000n V_low
+ 316.700001n V_low
+ 316.800000n V_low
+ 316.800001n V_low
+ 316.900000n V_low
+ 316.900001n V_low
+ 317.000000n V_low
+ 317.000001n V_low
+ 317.100000n V_low
+ 317.100001n V_low
+ 317.200000n V_low
+ 317.200001n V_low
+ 317.300000n V_low
+ 317.300001n V_low
+ 317.400000n V_low
+ 317.400001n V_low
+ 317.500000n V_low
+ 317.500001n V_low
+ 317.600000n V_low
+ 317.600001n V_low
+ 317.700000n V_low
+ 317.700001n V_low
+ 317.800000n V_low
+ 317.800001n V_low
+ 317.900000n V_low
+ 317.900001n V_low
+ 318.000000n V_low
+ 318.000001n V_hig
+ 318.100000n V_hig
+ 318.100001n V_hig
+ 318.200000n V_hig
+ 318.200001n V_hig
+ 318.300000n V_hig
+ 318.300001n V_hig
+ 318.400000n V_hig
+ 318.400001n V_hig
+ 318.500000n V_hig
+ 318.500001n V_hig
+ 318.600000n V_hig
+ 318.600001n V_hig
+ 318.700000n V_hig
+ 318.700001n V_hig
+ 318.800000n V_hig
+ 318.800001n V_hig
+ 318.900000n V_hig
+ 318.900001n V_hig
+ 319.000000n V_hig
+ 319.000001n V_hig
+ 319.100000n V_hig
+ 319.100001n V_hig
+ 319.200000n V_hig
+ 319.200001n V_hig
+ 319.300000n V_hig
+ 319.300001n V_hig
+ 319.400000n V_hig
+ 319.400001n V_hig
+ 319.500000n V_hig
+ 319.500001n V_hig
+ 319.600000n V_hig
+ 319.600001n V_hig
+ 319.700000n V_hig
+ 319.700001n V_hig
+ 319.800000n V_hig
+ 319.800001n V_hig
+ 319.900000n V_hig
+ 319.900001n V_hig
+ 320.000000n V_hig
+ 320.000001n V_hig
+ 320.100000n V_hig
+ 320.100001n V_hig
+ 320.200000n V_hig
+ 320.200001n V_hig
+ 320.300000n V_hig
+ 320.300001n V_hig
+ 320.400000n V_hig
+ 320.400001n V_hig
+ 320.500000n V_hig
+ 320.500001n V_hig
+ 320.600000n V_hig
+ 320.600001n V_hig
+ 320.700000n V_hig
+ 320.700001n V_hig
+ 320.800000n V_hig
+ 320.800001n V_hig
+ 320.900000n V_hig
+ 320.900001n V_hig
+ 321.000000n V_hig
+ 321.000001n V_low
+ 321.100000n V_low
+ 321.100001n V_low
+ 321.200000n V_low
+ 321.200001n V_low
+ 321.300000n V_low
+ 321.300001n V_low
+ 321.400000n V_low
+ 321.400001n V_low
+ 321.500000n V_low
+ 321.500001n V_low
+ 321.600000n V_low
+ 321.600001n V_low
+ 321.700000n V_low
+ 321.700001n V_low
+ 321.800000n V_low
+ 321.800001n V_low
+ 321.900000n V_low
+ 321.900001n V_low
+ 322.000000n V_low
+ 322.000001n V_low
+ 322.100000n V_low
+ 322.100001n V_low
+ 322.200000n V_low
+ 322.200001n V_low
+ 322.300000n V_low
+ 322.300001n V_low
+ 322.400000n V_low
+ 322.400001n V_low
+ 322.500000n V_low
+ 322.500001n V_low
+ 322.600000n V_low
+ 322.600001n V_low
+ 322.700000n V_low
+ 322.700001n V_low
+ 322.800000n V_low
+ 322.800001n V_low
+ 322.900000n V_low
+ 322.900001n V_low
+ 323.000000n V_low
+ 323.000001n V_low
+ 323.100000n V_low
+ 323.100001n V_low
+ 323.200000n V_low
+ 323.200001n V_low
+ 323.300000n V_low
+ 323.300001n V_low
+ 323.400000n V_low
+ 323.400001n V_low
+ 323.500000n V_low
+ 323.500001n V_low
+ 323.600000n V_low
+ 323.600001n V_low
+ 323.700000n V_low
+ 323.700001n V_low
+ 323.800000n V_low
+ 323.800001n V_low
+ 323.900000n V_low
+ 323.900001n V_low
+ 324.000000n V_low
+ 324.000001n V_hig
+ 324.100000n V_hig
+ 324.100001n V_hig
+ 324.200000n V_hig
+ 324.200001n V_hig
+ 324.300000n V_hig
+ 324.300001n V_hig
+ 324.400000n V_hig
+ 324.400001n V_hig
+ 324.500000n V_hig
+ 324.500001n V_hig
+ 324.600000n V_hig
+ 324.600001n V_hig
+ 324.700000n V_hig
+ 324.700001n V_hig
+ 324.800000n V_hig
+ 324.800001n V_hig
+ 324.900000n V_hig
+ 324.900001n V_hig
+ 325.000000n V_hig
+ 325.000001n V_hig
+ 325.100000n V_hig
+ 325.100001n V_hig
+ 325.200000n V_hig
+ 325.200001n V_hig
+ 325.300000n V_hig
+ 325.300001n V_hig
+ 325.400000n V_hig
+ 325.400001n V_hig
+ 325.500000n V_hig
+ 325.500001n V_hig
+ 325.600000n V_hig
+ 325.600001n V_hig
+ 325.700000n V_hig
+ 325.700001n V_hig
+ 325.800000n V_hig
+ 325.800001n V_hig
+ 325.900000n V_hig
+ 325.900001n V_hig
+ 326.000000n V_hig
+ 326.000001n V_low
+ 326.100000n V_low
+ 326.100001n V_low
+ 326.200000n V_low
+ 326.200001n V_low
+ 326.300000n V_low
+ 326.300001n V_low
+ 326.400000n V_low
+ 326.400001n V_low
+ 326.500000n V_low
+ 326.500001n V_low
+ 326.600000n V_low
+ 326.600001n V_low
+ 326.700000n V_low
+ 326.700001n V_low
+ 326.800000n V_low
+ 326.800001n V_low
+ 326.900000n V_low
+ 326.900001n V_low
+ 327.000000n V_low
+ 327.000001n V_hig
+ 327.100000n V_hig
+ 327.100001n V_hig
+ 327.200000n V_hig
+ 327.200001n V_hig
+ 327.300000n V_hig
+ 327.300001n V_hig
+ 327.400000n V_hig
+ 327.400001n V_hig
+ 327.500000n V_hig
+ 327.500001n V_hig
+ 327.600000n V_hig
+ 327.600001n V_hig
+ 327.700000n V_hig
+ 327.700001n V_hig
+ 327.800000n V_hig
+ 327.800001n V_hig
+ 327.900000n V_hig
+ 327.900001n V_hig
+ 328.000000n V_hig
+ 328.000001n V_low
+ 328.100000n V_low
+ 328.100001n V_low
+ 328.200000n V_low
+ 328.200001n V_low
+ 328.300000n V_low
+ 328.300001n V_low
+ 328.400000n V_low
+ 328.400001n V_low
+ 328.500000n V_low
+ 328.500001n V_low
+ 328.600000n V_low
+ 328.600001n V_low
+ 328.700000n V_low
+ 328.700001n V_low
+ 328.800000n V_low
+ 328.800001n V_low
+ 328.900000n V_low
+ 328.900001n V_low
+ 329.000000n V_low
+ 329.000001n V_hig
+ 329.100000n V_hig
+ 329.100001n V_hig
+ 329.200000n V_hig
+ 329.200001n V_hig
+ 329.300000n V_hig
+ 329.300001n V_hig
+ 329.400000n V_hig
+ 329.400001n V_hig
+ 329.500000n V_hig
+ 329.500001n V_hig
+ 329.600000n V_hig
+ 329.600001n V_hig
+ 329.700000n V_hig
+ 329.700001n V_hig
+ 329.800000n V_hig
+ 329.800001n V_hig
+ 329.900000n V_hig
+ 329.900001n V_hig
+ 330.000000n V_hig
+ 330.000001n V_low
+ 330.100000n V_low
+ 330.100001n V_low
+ 330.200000n V_low
+ 330.200001n V_low
+ 330.300000n V_low
+ 330.300001n V_low
+ 330.400000n V_low
+ 330.400001n V_low
+ 330.500000n V_low
+ 330.500001n V_low
+ 330.600000n V_low
+ 330.600001n V_low
+ 330.700000n V_low
+ 330.700001n V_low
+ 330.800000n V_low
+ 330.800001n V_low
+ 330.900000n V_low
+ 330.900001n V_low
+ 331.000000n V_low
+ 331.000001n V_low
+ 331.100000n V_low
+ 331.100001n V_low
+ 331.200000n V_low
+ 331.200001n V_low
+ 331.300000n V_low
+ 331.300001n V_low
+ 331.400000n V_low
+ 331.400001n V_low
+ 331.500000n V_low
+ 331.500001n V_low
+ 331.600000n V_low
+ 331.600001n V_low
+ 331.700000n V_low
+ 331.700001n V_low
+ 331.800000n V_low
+ 331.800001n V_low
+ 331.900000n V_low
+ 331.900001n V_low
+ 332.000000n V_low
+ 332.000001n V_hig
+ 332.100000n V_hig
+ 332.100001n V_hig
+ 332.200000n V_hig
+ 332.200001n V_hig
+ 332.300000n V_hig
+ 332.300001n V_hig
+ 332.400000n V_hig
+ 332.400001n V_hig
+ 332.500000n V_hig
+ 332.500001n V_hig
+ 332.600000n V_hig
+ 332.600001n V_hig
+ 332.700000n V_hig
+ 332.700001n V_hig
+ 332.800000n V_hig
+ 332.800001n V_hig
+ 332.900000n V_hig
+ 332.900001n V_hig
+ 333.000000n V_hig
+ 333.000001n V_hig
+ 333.100000n V_hig
+ 333.100001n V_hig
+ 333.200000n V_hig
+ 333.200001n V_hig
+ 333.300000n V_hig
+ 333.300001n V_hig
+ 333.400000n V_hig
+ 333.400001n V_hig
+ 333.500000n V_hig
+ 333.500001n V_hig
+ 333.600000n V_hig
+ 333.600001n V_hig
+ 333.700000n V_hig
+ 333.700001n V_hig
+ 333.800000n V_hig
+ 333.800001n V_hig
+ 333.900000n V_hig
+ 333.900001n V_hig
+ 334.000000n V_hig
+ 334.000001n V_hig
+ 334.100000n V_hig
+ 334.100001n V_hig
+ 334.200000n V_hig
+ 334.200001n V_hig
+ 334.300000n V_hig
+ 334.300001n V_hig
+ 334.400000n V_hig
+ 334.400001n V_hig
+ 334.500000n V_hig
+ 334.500001n V_hig
+ 334.600000n V_hig
+ 334.600001n V_hig
+ 334.700000n V_hig
+ 334.700001n V_hig
+ 334.800000n V_hig
+ 334.800001n V_hig
+ 334.900000n V_hig
+ 334.900001n V_hig
+ 335.000000n V_hig
+ 335.000001n V_hig
+ 335.100000n V_hig
+ 335.100001n V_hig
+ 335.200000n V_hig
+ 335.200001n V_hig
+ 335.300000n V_hig
+ 335.300001n V_hig
+ 335.400000n V_hig
+ 335.400001n V_hig
+ 335.500000n V_hig
+ 335.500001n V_hig
+ 335.600000n V_hig
+ 335.600001n V_hig
+ 335.700000n V_hig
+ 335.700001n V_hig
+ 335.800000n V_hig
+ 335.800001n V_hig
+ 335.900000n V_hig
+ 335.900001n V_hig
+ 336.000000n V_hig
+ 336.000001n V_low
+ 336.100000n V_low
+ 336.100001n V_low
+ 336.200000n V_low
+ 336.200001n V_low
+ 336.300000n V_low
+ 336.300001n V_low
+ 336.400000n V_low
+ 336.400001n V_low
+ 336.500000n V_low
+ 336.500001n V_low
+ 336.600000n V_low
+ 336.600001n V_low
+ 336.700000n V_low
+ 336.700001n V_low
+ 336.800000n V_low
+ 336.800001n V_low
+ 336.900000n V_low
+ 336.900001n V_low
+ 337.000000n V_low
+ 337.000001n V_hig
+ 337.100000n V_hig
+ 337.100001n V_hig
+ 337.200000n V_hig
+ 337.200001n V_hig
+ 337.300000n V_hig
+ 337.300001n V_hig
+ 337.400000n V_hig
+ 337.400001n V_hig
+ 337.500000n V_hig
+ 337.500001n V_hig
+ 337.600000n V_hig
+ 337.600001n V_hig
+ 337.700000n V_hig
+ 337.700001n V_hig
+ 337.800000n V_hig
+ 337.800001n V_hig
+ 337.900000n V_hig
+ 337.900001n V_hig
+ 338.000000n V_hig
+ 338.000001n V_low
+ 338.100000n V_low
+ 338.100001n V_low
+ 338.200000n V_low
+ 338.200001n V_low
+ 338.300000n V_low
+ 338.300001n V_low
+ 338.400000n V_low
+ 338.400001n V_low
+ 338.500000n V_low
+ 338.500001n V_low
+ 338.600000n V_low
+ 338.600001n V_low
+ 338.700000n V_low
+ 338.700001n V_low
+ 338.800000n V_low
+ 338.800001n V_low
+ 338.900000n V_low
+ 338.900001n V_low
+ 339.000000n V_low
+ 339.000001n V_low
+ 339.100000n V_low
+ 339.100001n V_low
+ 339.200000n V_low
+ 339.200001n V_low
+ 339.300000n V_low
+ 339.300001n V_low
+ 339.400000n V_low
+ 339.400001n V_low
+ 339.500000n V_low
+ 339.500001n V_low
+ 339.600000n V_low
+ 339.600001n V_low
+ 339.700000n V_low
+ 339.700001n V_low
+ 339.800000n V_low
+ 339.800001n V_low
+ 339.900000n V_low
+ 339.900001n V_low
+ 340.000000n V_low
+ 340.000001n V_low
+ 340.100000n V_low
+ 340.100001n V_low
+ 340.200000n V_low
+ 340.200001n V_low
+ 340.300000n V_low
+ 340.300001n V_low
+ 340.400000n V_low
+ 340.400001n V_low
+ 340.500000n V_low
+ 340.500001n V_low
+ 340.600000n V_low
+ 340.600001n V_low
+ 340.700000n V_low
+ 340.700001n V_low
+ 340.800000n V_low
+ 340.800001n V_low
+ 340.900000n V_low
+ 340.900001n V_low
+ 341.000000n V_low
+ 341.000001n V_hig
+ 341.100000n V_hig
+ 341.100001n V_hig
+ 341.200000n V_hig
+ 341.200001n V_hig
+ 341.300000n V_hig
+ 341.300001n V_hig
+ 341.400000n V_hig
+ 341.400001n V_hig
+ 341.500000n V_hig
+ 341.500001n V_hig
+ 341.600000n V_hig
+ 341.600001n V_hig
+ 341.700000n V_hig
+ 341.700001n V_hig
+ 341.800000n V_hig
+ 341.800001n V_hig
+ 341.900000n V_hig
+ 341.900001n V_hig
+ 342.000000n V_hig
+ 342.000001n V_hig
+ 342.100000n V_hig
+ 342.100001n V_hig
+ 342.200000n V_hig
+ 342.200001n V_hig
+ 342.300000n V_hig
+ 342.300001n V_hig
+ 342.400000n V_hig
+ 342.400001n V_hig
+ 342.500000n V_hig
+ 342.500001n V_hig
+ 342.600000n V_hig
+ 342.600001n V_hig
+ 342.700000n V_hig
+ 342.700001n V_hig
+ 342.800000n V_hig
+ 342.800001n V_hig
+ 342.900000n V_hig
+ 342.900001n V_hig
+ 343.000000n V_hig
+ 343.000001n V_low
+ 343.100000n V_low
+ 343.100001n V_low
+ 343.200000n V_low
+ 343.200001n V_low
+ 343.300000n V_low
+ 343.300001n V_low
+ 343.400000n V_low
+ 343.400001n V_low
+ 343.500000n V_low
+ 343.500001n V_low
+ 343.600000n V_low
+ 343.600001n V_low
+ 343.700000n V_low
+ 343.700001n V_low
+ 343.800000n V_low
+ 343.800001n V_low
+ 343.900000n V_low
+ 343.900001n V_low
+ 344.000000n V_low
+ 344.000001n V_hig
+ 344.100000n V_hig
+ 344.100001n V_hig
+ 344.200000n V_hig
+ 344.200001n V_hig
+ 344.300000n V_hig
+ 344.300001n V_hig
+ 344.400000n V_hig
+ 344.400001n V_hig
+ 344.500000n V_hig
+ 344.500001n V_hig
+ 344.600000n V_hig
+ 344.600001n V_hig
+ 344.700000n V_hig
+ 344.700001n V_hig
+ 344.800000n V_hig
+ 344.800001n V_hig
+ 344.900000n V_hig
+ 344.900001n V_hig
+ 345.000000n V_hig
+ 345.000001n V_hig
+ 345.100000n V_hig
+ 345.100001n V_hig
+ 345.200000n V_hig
+ 345.200001n V_hig
+ 345.300000n V_hig
+ 345.300001n V_hig
+ 345.400000n V_hig
+ 345.400001n V_hig
+ 345.500000n V_hig
+ 345.500001n V_hig
+ 345.600000n V_hig
+ 345.600001n V_hig
+ 345.700000n V_hig
+ 345.700001n V_hig
+ 345.800000n V_hig
+ 345.800001n V_hig
+ 345.900000n V_hig
+ 345.900001n V_hig
+ 346.000000n V_hig
+ 346.000001n V_low
+ 346.100000n V_low
+ 346.100001n V_low
+ 346.200000n V_low
+ 346.200001n V_low
+ 346.300000n V_low
+ 346.300001n V_low
+ 346.400000n V_low
+ 346.400001n V_low
+ 346.500000n V_low
+ 346.500001n V_low
+ 346.600000n V_low
+ 346.600001n V_low
+ 346.700000n V_low
+ 346.700001n V_low
+ 346.800000n V_low
+ 346.800001n V_low
+ 346.900000n V_low
+ 346.900001n V_low
+ 347.000000n V_low
+ 347.000001n V_low
+ 347.100000n V_low
+ 347.100001n V_low
+ 347.200000n V_low
+ 347.200001n V_low
+ 347.300000n V_low
+ 347.300001n V_low
+ 347.400000n V_low
+ 347.400001n V_low
+ 347.500000n V_low
+ 347.500001n V_low
+ 347.600000n V_low
+ 347.600001n V_low
+ 347.700000n V_low
+ 347.700001n V_low
+ 347.800000n V_low
+ 347.800001n V_low
+ 347.900000n V_low
+ 347.900001n V_low
+ 348.000000n V_low
+ 348.000001n V_low
+ 348.100000n V_low
+ 348.100001n V_low
+ 348.200000n V_low
+ 348.200001n V_low
+ 348.300000n V_low
+ 348.300001n V_low
+ 348.400000n V_low
+ 348.400001n V_low
+ 348.500000n V_low
+ 348.500001n V_low
+ 348.600000n V_low
+ 348.600001n V_low
+ 348.700000n V_low
+ 348.700001n V_low
+ 348.800000n V_low
+ 348.800001n V_low
+ 348.900000n V_low
+ 348.900001n V_low
+ 349.000000n V_low
+ 349.000001n V_hig
+ 349.100000n V_hig
+ 349.100001n V_hig
+ 349.200000n V_hig
+ 349.200001n V_hig
+ 349.300000n V_hig
+ 349.300001n V_hig
+ 349.400000n V_hig
+ 349.400001n V_hig
+ 349.500000n V_hig
+ 349.500001n V_hig
+ 349.600000n V_hig
+ 349.600001n V_hig
+ 349.700000n V_hig
+ 349.700001n V_hig
+ 349.800000n V_hig
+ 349.800001n V_hig
+ 349.900000n V_hig
+ 349.900001n V_hig
+ 350.000000n V_hig
+ 350.000001n V_hig
+ 350.100000n V_hig
+ 350.100001n V_hig
+ 350.200000n V_hig
+ 350.200001n V_hig
+ 350.300000n V_hig
+ 350.300001n V_hig
+ 350.400000n V_hig
+ 350.400001n V_hig
+ 350.500000n V_hig
+ 350.500001n V_hig
+ 350.600000n V_hig
+ 350.600001n V_hig
+ 350.700000n V_hig
+ 350.700001n V_hig
+ 350.800000n V_hig
+ 350.800001n V_hig
+ 350.900000n V_hig
+ 350.900001n V_hig
+ 351.000000n V_hig
+ 351.000001n V_hig
+ 351.100000n V_hig
+ 351.100001n V_hig
+ 351.200000n V_hig
+ 351.200001n V_hig
+ 351.300000n V_hig
+ 351.300001n V_hig
+ 351.400000n V_hig
+ 351.400001n V_hig
+ 351.500000n V_hig
+ 351.500001n V_hig
+ 351.600000n V_hig
+ 351.600001n V_hig
+ 351.700000n V_hig
+ 351.700001n V_hig
+ 351.800000n V_hig
+ 351.800001n V_hig
+ 351.900000n V_hig
+ 351.900001n V_hig
+ 352.000000n V_hig
+ 352.000001n V_hig
+ 352.100000n V_hig
+ 352.100001n V_hig
+ 352.200000n V_hig
+ 352.200001n V_hig
+ 352.300000n V_hig
+ 352.300001n V_hig
+ 352.400000n V_hig
+ 352.400001n V_hig
+ 352.500000n V_hig
+ 352.500001n V_hig
+ 352.600000n V_hig
+ 352.600001n V_hig
+ 352.700000n V_hig
+ 352.700001n V_hig
+ 352.800000n V_hig
+ 352.800001n V_hig
+ 352.900000n V_hig
+ 352.900001n V_hig
+ 353.000000n V_hig
+ 353.000001n V_hig
+ 353.100000n V_hig
+ 353.100001n V_hig
+ 353.200000n V_hig
+ 353.200001n V_hig
+ 353.300000n V_hig
+ 353.300001n V_hig
+ 353.400000n V_hig
+ 353.400001n V_hig
+ 353.500000n V_hig
+ 353.500001n V_hig
+ 353.600000n V_hig
+ 353.600001n V_hig
+ 353.700000n V_hig
+ 353.700001n V_hig
+ 353.800000n V_hig
+ 353.800001n V_hig
+ 353.900000n V_hig
+ 353.900001n V_hig
+ 354.000000n V_hig
+ 354.000001n V_hig
+ 354.100000n V_hig
+ 354.100001n V_hig
+ 354.200000n V_hig
+ 354.200001n V_hig
+ 354.300000n V_hig
+ 354.300001n V_hig
+ 354.400000n V_hig
+ 354.400001n V_hig
+ 354.500000n V_hig
+ 354.500001n V_hig
+ 354.600000n V_hig
+ 354.600001n V_hig
+ 354.700000n V_hig
+ 354.700001n V_hig
+ 354.800000n V_hig
+ 354.800001n V_hig
+ 354.900000n V_hig
+ 354.900001n V_hig
+ 355.000000n V_hig
+ 355.000001n V_hig
+ 355.100000n V_hig
+ 355.100001n V_hig
+ 355.200000n V_hig
+ 355.200001n V_hig
+ 355.300000n V_hig
+ 355.300001n V_hig
+ 355.400000n V_hig
+ 355.400001n V_hig
+ 355.500000n V_hig
+ 355.500001n V_hig
+ 355.600000n V_hig
+ 355.600001n V_hig
+ 355.700000n V_hig
+ 355.700001n V_hig
+ 355.800000n V_hig
+ 355.800001n V_hig
+ 355.900000n V_hig
+ 355.900001n V_hig
+ 356.000000n V_hig
+ 356.000001n V_hig
+ 356.100000n V_hig
+ 356.100001n V_hig
+ 356.200000n V_hig
+ 356.200001n V_hig
+ 356.300000n V_hig
+ 356.300001n V_hig
+ 356.400000n V_hig
+ 356.400001n V_hig
+ 356.500000n V_hig
+ 356.500001n V_hig
+ 356.600000n V_hig
+ 356.600001n V_hig
+ 356.700000n V_hig
+ 356.700001n V_hig
+ 356.800000n V_hig
+ 356.800001n V_hig
+ 356.900000n V_hig
+ 356.900001n V_hig
+ 357.000000n V_hig
+ 357.000001n V_low
+ 357.100000n V_low
+ 357.100001n V_low
+ 357.200000n V_low
+ 357.200001n V_low
+ 357.300000n V_low
+ 357.300001n V_low
+ 357.400000n V_low
+ 357.400001n V_low
+ 357.500000n V_low
+ 357.500001n V_low
+ 357.600000n V_low
+ 357.600001n V_low
+ 357.700000n V_low
+ 357.700001n V_low
+ 357.800000n V_low
+ 357.800001n V_low
+ 357.900000n V_low
+ 357.900001n V_low
+ 358.000000n V_low
+ 358.000001n V_hig
+ 358.100000n V_hig
+ 358.100001n V_hig
+ 358.200000n V_hig
+ 358.200001n V_hig
+ 358.300000n V_hig
+ 358.300001n V_hig
+ 358.400000n V_hig
+ 358.400001n V_hig
+ 358.500000n V_hig
+ 358.500001n V_hig
+ 358.600000n V_hig
+ 358.600001n V_hig
+ 358.700000n V_hig
+ 358.700001n V_hig
+ 358.800000n V_hig
+ 358.800001n V_hig
+ 358.900000n V_hig
+ 358.900001n V_hig
+ 359.000000n V_hig
+ 359.000001n V_low
+ 359.100000n V_low
+ 359.100001n V_low
+ 359.200000n V_low
+ 359.200001n V_low
+ 359.300000n V_low
+ 359.300001n V_low
+ 359.400000n V_low
+ 359.400001n V_low
+ 359.500000n V_low
+ 359.500001n V_low
+ 359.600000n V_low
+ 359.600001n V_low
+ 359.700000n V_low
+ 359.700001n V_low
+ 359.800000n V_low
+ 359.800001n V_low
+ 359.900000n V_low
+ 359.900001n V_low
+ 360.000000n V_low
+ 360.000001n V_hig
+ 360.100000n V_hig
+ 360.100001n V_hig
+ 360.200000n V_hig
+ 360.200001n V_hig
+ 360.300000n V_hig
+ 360.300001n V_hig
+ 360.400000n V_hig
+ 360.400001n V_hig
+ 360.500000n V_hig
+ 360.500001n V_hig
+ 360.600000n V_hig
+ 360.600001n V_hig
+ 360.700000n V_hig
+ 360.700001n V_hig
+ 360.800000n V_hig
+ 360.800001n V_hig
+ 360.900000n V_hig
+ 360.900001n V_hig
+ 361.000000n V_hig
+ 361.000001n V_hig
+ 361.100000n V_hig
+ 361.100001n V_hig
+ 361.200000n V_hig
+ 361.200001n V_hig
+ 361.300000n V_hig
+ 361.300001n V_hig
+ 361.400000n V_hig
+ 361.400001n V_hig
+ 361.500000n V_hig
+ 361.500001n V_hig
+ 361.600000n V_hig
+ 361.600001n V_hig
+ 361.700000n V_hig
+ 361.700001n V_hig
+ 361.800000n V_hig
+ 361.800001n V_hig
+ 361.900000n V_hig
+ 361.900001n V_hig
+ 362.000000n V_hig
+ 362.000001n V_hig
+ 362.100000n V_hig
+ 362.100001n V_hig
+ 362.200000n V_hig
+ 362.200001n V_hig
+ 362.300000n V_hig
+ 362.300001n V_hig
+ 362.400000n V_hig
+ 362.400001n V_hig
+ 362.500000n V_hig
+ 362.500001n V_hig
+ 362.600000n V_hig
+ 362.600001n V_hig
+ 362.700000n V_hig
+ 362.700001n V_hig
+ 362.800000n V_hig
+ 362.800001n V_hig
+ 362.900000n V_hig
+ 362.900001n V_hig
+ 363.000000n V_hig
+ 363.000001n V_low
+ 363.100000n V_low
+ 363.100001n V_low
+ 363.200000n V_low
+ 363.200001n V_low
+ 363.300000n V_low
+ 363.300001n V_low
+ 363.400000n V_low
+ 363.400001n V_low
+ 363.500000n V_low
+ 363.500001n V_low
+ 363.600000n V_low
+ 363.600001n V_low
+ 363.700000n V_low
+ 363.700001n V_low
+ 363.800000n V_low
+ 363.800001n V_low
+ 363.900000n V_low
+ 363.900001n V_low
+ 364.000000n V_low
+ 364.000001n V_hig
+ 364.100000n V_hig
+ 364.100001n V_hig
+ 364.200000n V_hig
+ 364.200001n V_hig
+ 364.300000n V_hig
+ 364.300001n V_hig
+ 364.400000n V_hig
+ 364.400001n V_hig
+ 364.500000n V_hig
+ 364.500001n V_hig
+ 364.600000n V_hig
+ 364.600001n V_hig
+ 364.700000n V_hig
+ 364.700001n V_hig
+ 364.800000n V_hig
+ 364.800001n V_hig
+ 364.900000n V_hig
+ 364.900001n V_hig
+ 365.000000n V_hig
+ 365.000001n V_low
+ 365.100000n V_low
+ 365.100001n V_low
+ 365.200000n V_low
+ 365.200001n V_low
+ 365.300000n V_low
+ 365.300001n V_low
+ 365.400000n V_low
+ 365.400001n V_low
+ 365.500000n V_low
+ 365.500001n V_low
+ 365.600000n V_low
+ 365.600001n V_low
+ 365.700000n V_low
+ 365.700001n V_low
+ 365.800000n V_low
+ 365.800001n V_low
+ 365.900000n V_low
+ 365.900001n V_low
+ 366.000000n V_low
+ 366.000001n V_hig
+ 366.100000n V_hig
+ 366.100001n V_hig
+ 366.200000n V_hig
+ 366.200001n V_hig
+ 366.300000n V_hig
+ 366.300001n V_hig
+ 366.400000n V_hig
+ 366.400001n V_hig
+ 366.500000n V_hig
+ 366.500001n V_hig
+ 366.600000n V_hig
+ 366.600001n V_hig
+ 366.700000n V_hig
+ 366.700001n V_hig
+ 366.800000n V_hig
+ 366.800001n V_hig
+ 366.900000n V_hig
+ 366.900001n V_hig
+ 367.000000n V_hig
+ 367.000001n V_hig
+ 367.100000n V_hig
+ 367.100001n V_hig
+ 367.200000n V_hig
+ 367.200001n V_hig
+ 367.300000n V_hig
+ 367.300001n V_hig
+ 367.400000n V_hig
+ 367.400001n V_hig
+ 367.500000n V_hig
+ 367.500001n V_hig
+ 367.600000n V_hig
+ 367.600001n V_hig
+ 367.700000n V_hig
+ 367.700001n V_hig
+ 367.800000n V_hig
+ 367.800001n V_hig
+ 367.900000n V_hig
+ 367.900001n V_hig
+ 368.000000n V_hig
+ 368.000001n V_low
+ 368.100000n V_low
+ 368.100001n V_low
+ 368.200000n V_low
+ 368.200001n V_low
+ 368.300000n V_low
+ 368.300001n V_low
+ 368.400000n V_low
+ 368.400001n V_low
+ 368.500000n V_low
+ 368.500001n V_low
+ 368.600000n V_low
+ 368.600001n V_low
+ 368.700000n V_low
+ 368.700001n V_low
+ 368.800000n V_low
+ 368.800001n V_low
+ 368.900000n V_low
+ 368.900001n V_low
+ 369.000000n V_low
+ 369.000001n V_hig
+ 369.100000n V_hig
+ 369.100001n V_hig
+ 369.200000n V_hig
+ 369.200001n V_hig
+ 369.300000n V_hig
+ 369.300001n V_hig
+ 369.400000n V_hig
+ 369.400001n V_hig
+ 369.500000n V_hig
+ 369.500001n V_hig
+ 369.600000n V_hig
+ 369.600001n V_hig
+ 369.700000n V_hig
+ 369.700001n V_hig
+ 369.800000n V_hig
+ 369.800001n V_hig
+ 369.900000n V_hig
+ 369.900001n V_hig
+ 370.000000n V_hig
+ 370.000001n V_low
+ 370.100000n V_low
+ 370.100001n V_low
+ 370.200000n V_low
+ 370.200001n V_low
+ 370.300000n V_low
+ 370.300001n V_low
+ 370.400000n V_low
+ 370.400001n V_low
+ 370.500000n V_low
+ 370.500001n V_low
+ 370.600000n V_low
+ 370.600001n V_low
+ 370.700000n V_low
+ 370.700001n V_low
+ 370.800000n V_low
+ 370.800001n V_low
+ 370.900000n V_low
+ 370.900001n V_low
+ 371.000000n V_low
+ 371.000001n V_hig
+ 371.100000n V_hig
+ 371.100001n V_hig
+ 371.200000n V_hig
+ 371.200001n V_hig
+ 371.300000n V_hig
+ 371.300001n V_hig
+ 371.400000n V_hig
+ 371.400001n V_hig
+ 371.500000n V_hig
+ 371.500001n V_hig
+ 371.600000n V_hig
+ 371.600001n V_hig
+ 371.700000n V_hig
+ 371.700001n V_hig
+ 371.800000n V_hig
+ 371.800001n V_hig
+ 371.900000n V_hig
+ 371.900001n V_hig
+ 372.000000n V_hig
+ 372.000001n V_low
+ 372.100000n V_low
+ 372.100001n V_low
+ 372.200000n V_low
+ 372.200001n V_low
+ 372.300000n V_low
+ 372.300001n V_low
+ 372.400000n V_low
+ 372.400001n V_low
+ 372.500000n V_low
+ 372.500001n V_low
+ 372.600000n V_low
+ 372.600001n V_low
+ 372.700000n V_low
+ 372.700001n V_low
+ 372.800000n V_low
+ 372.800001n V_low
+ 372.900000n V_low
+ 372.900001n V_low
+ 373.000000n V_low
+ 373.000001n V_hig
+ 373.100000n V_hig
+ 373.100001n V_hig
+ 373.200000n V_hig
+ 373.200001n V_hig
+ 373.300000n V_hig
+ 373.300001n V_hig
+ 373.400000n V_hig
+ 373.400001n V_hig
+ 373.500000n V_hig
+ 373.500001n V_hig
+ 373.600000n V_hig
+ 373.600001n V_hig
+ 373.700000n V_hig
+ 373.700001n V_hig
+ 373.800000n V_hig
+ 373.800001n V_hig
+ 373.900000n V_hig
+ 373.900001n V_hig
+ 374.000000n V_hig
+ 374.000001n V_hig
+ 374.100000n V_hig
+ 374.100001n V_hig
+ 374.200000n V_hig
+ 374.200001n V_hig
+ 374.300000n V_hig
+ 374.300001n V_hig
+ 374.400000n V_hig
+ 374.400001n V_hig
+ 374.500000n V_hig
+ 374.500001n V_hig
+ 374.600000n V_hig
+ 374.600001n V_hig
+ 374.700000n V_hig
+ 374.700001n V_hig
+ 374.800000n V_hig
+ 374.800001n V_hig
+ 374.900000n V_hig
+ 374.900001n V_hig
+ 375.000000n V_hig
+ 375.000001n V_hig
+ 375.100000n V_hig
+ 375.100001n V_hig
+ 375.200000n V_hig
+ 375.200001n V_hig
+ 375.300000n V_hig
+ 375.300001n V_hig
+ 375.400000n V_hig
+ 375.400001n V_hig
+ 375.500000n V_hig
+ 375.500001n V_hig
+ 375.600000n V_hig
+ 375.600001n V_hig
+ 375.700000n V_hig
+ 375.700001n V_hig
+ 375.800000n V_hig
+ 375.800001n V_hig
+ 375.900000n V_hig
+ 375.900001n V_hig
+ 376.000000n V_hig
+ 376.000001n V_hig
+ 376.100000n V_hig
+ 376.100001n V_hig
+ 376.200000n V_hig
+ 376.200001n V_hig
+ 376.300000n V_hig
+ 376.300001n V_hig
+ 376.400000n V_hig
+ 376.400001n V_hig
+ 376.500000n V_hig
+ 376.500001n V_hig
+ 376.600000n V_hig
+ 376.600001n V_hig
+ 376.700000n V_hig
+ 376.700001n V_hig
+ 376.800000n V_hig
+ 376.800001n V_hig
+ 376.900000n V_hig
+ 376.900001n V_hig
+ 377.000000n V_hig
+ 377.000001n V_low
+ 377.100000n V_low
+ 377.100001n V_low
+ 377.200000n V_low
+ 377.200001n V_low
+ 377.300000n V_low
+ 377.300001n V_low
+ 377.400000n V_low
+ 377.400001n V_low
+ 377.500000n V_low
+ 377.500001n V_low
+ 377.600000n V_low
+ 377.600001n V_low
+ 377.700000n V_low
+ 377.700001n V_low
+ 377.800000n V_low
+ 377.800001n V_low
+ 377.900000n V_low
+ 377.900001n V_low
+ 378.000000n V_low
+ 378.000001n V_low
+ 378.100000n V_low
+ 378.100001n V_low
+ 378.200000n V_low
+ 378.200001n V_low
+ 378.300000n V_low
+ 378.300001n V_low
+ 378.400000n V_low
+ 378.400001n V_low
+ 378.500000n V_low
+ 378.500001n V_low
+ 378.600000n V_low
+ 378.600001n V_low
+ 378.700000n V_low
+ 378.700001n V_low
+ 378.800000n V_low
+ 378.800001n V_low
+ 378.900000n V_low
+ 378.900001n V_low
+ 379.000000n V_low
+ 379.000001n V_low
+ 379.100000n V_low
+ 379.100001n V_low
+ 379.200000n V_low
+ 379.200001n V_low
+ 379.300000n V_low
+ 379.300001n V_low
+ 379.400000n V_low
+ 379.400001n V_low
+ 379.500000n V_low
+ 379.500001n V_low
+ 379.600000n V_low
+ 379.600001n V_low
+ 379.700000n V_low
+ 379.700001n V_low
+ 379.800000n V_low
+ 379.800001n V_low
+ 379.900000n V_low
+ 379.900001n V_low
+ 380.000000n V_low
+ 380.000001n V_low
+ 380.100000n V_low
+ 380.100001n V_low
+ 380.200000n V_low
+ 380.200001n V_low
+ 380.300000n V_low
+ 380.300001n V_low
+ 380.400000n V_low
+ 380.400001n V_low
+ 380.500000n V_low
+ 380.500001n V_low
+ 380.600000n V_low
+ 380.600001n V_low
+ 380.700000n V_low
+ 380.700001n V_low
+ 380.800000n V_low
+ 380.800001n V_low
+ 380.900000n V_low
+ 380.900001n V_low
+ 381.000000n V_low
+ 381.000001n V_hig
+ 381.100000n V_hig
+ 381.100001n V_hig
+ 381.200000n V_hig
+ 381.200001n V_hig
+ 381.300000n V_hig
+ 381.300001n V_hig
+ 381.400000n V_hig
+ 381.400001n V_hig
+ 381.500000n V_hig
+ 381.500001n V_hig
+ 381.600000n V_hig
+ 381.600001n V_hig
+ 381.700000n V_hig
+ 381.700001n V_hig
+ 381.800000n V_hig
+ 381.800001n V_hig
+ 381.900000n V_hig
+ 381.900001n V_hig
+ 382.000000n V_hig
+ 382.000001n V_hig
+ 382.100000n V_hig
+ 382.100001n V_hig
+ 382.200000n V_hig
+ 382.200001n V_hig
+ 382.300000n V_hig
+ 382.300001n V_hig
+ 382.400000n V_hig
+ 382.400001n V_hig
+ 382.500000n V_hig
+ 382.500001n V_hig
+ 382.600000n V_hig
+ 382.600001n V_hig
+ 382.700000n V_hig
+ 382.700001n V_hig
+ 382.800000n V_hig
+ 382.800001n V_hig
+ 382.900000n V_hig
+ 382.900001n V_hig
+ 383.000000n V_hig
+ 383.000001n V_low
+ 383.100000n V_low
+ 383.100001n V_low
+ 383.200000n V_low
+ 383.200001n V_low
+ 383.300000n V_low
+ 383.300001n V_low
+ 383.400000n V_low
+ 383.400001n V_low
+ 383.500000n V_low
+ 383.500001n V_low
+ 383.600000n V_low
+ 383.600001n V_low
+ 383.700000n V_low
+ 383.700001n V_low
+ 383.800000n V_low
+ 383.800001n V_low
+ 383.900000n V_low
+ 383.900001n V_low
+ 384.000000n V_low
+ 384.000001n V_hig
+ 384.100000n V_hig
+ 384.100001n V_hig
+ 384.200000n V_hig
+ 384.200001n V_hig
+ 384.300000n V_hig
+ 384.300001n V_hig
+ 384.400000n V_hig
+ 384.400001n V_hig
+ 384.500000n V_hig
+ 384.500001n V_hig
+ 384.600000n V_hig
+ 384.600001n V_hig
+ 384.700000n V_hig
+ 384.700001n V_hig
+ 384.800000n V_hig
+ 384.800001n V_hig
+ 384.900000n V_hig
+ 384.900001n V_hig
+ 385.000000n V_hig
+ 385.000001n V_low
+ 385.100000n V_low
+ 385.100001n V_low
+ 385.200000n V_low
+ 385.200001n V_low
+ 385.300000n V_low
+ 385.300001n V_low
+ 385.400000n V_low
+ 385.400001n V_low
+ 385.500000n V_low
+ 385.500001n V_low
+ 385.600000n V_low
+ 385.600001n V_low
+ 385.700000n V_low
+ 385.700001n V_low
+ 385.800000n V_low
+ 385.800001n V_low
+ 385.900000n V_low
+ 385.900001n V_low
+ 386.000000n V_low
+ 386.000001n V_low
+ 386.100000n V_low
+ 386.100001n V_low
+ 386.200000n V_low
+ 386.200001n V_low
+ 386.300000n V_low
+ 386.300001n V_low
+ 386.400000n V_low
+ 386.400001n V_low
+ 386.500000n V_low
+ 386.500001n V_low
+ 386.600000n V_low
+ 386.600001n V_low
+ 386.700000n V_low
+ 386.700001n V_low
+ 386.800000n V_low
+ 386.800001n V_low
+ 386.900000n V_low
+ 386.900001n V_low
+ 387.000000n V_low
+ 387.000001n V_low
+ 387.100000n V_low
+ 387.100001n V_low
+ 387.200000n V_low
+ 387.200001n V_low
+ 387.300000n V_low
+ 387.300001n V_low
+ 387.400000n V_low
+ 387.400001n V_low
+ 387.500000n V_low
+ 387.500001n V_low
+ 387.600000n V_low
+ 387.600001n V_low
+ 387.700000n V_low
+ 387.700001n V_low
+ 387.800000n V_low
+ 387.800001n V_low
+ 387.900000n V_low
+ 387.900001n V_low
+ 388.000000n V_low
+ 388.000001n V_hig
+ 388.100000n V_hig
+ 388.100001n V_hig
+ 388.200000n V_hig
+ 388.200001n V_hig
+ 388.300000n V_hig
+ 388.300001n V_hig
+ 388.400000n V_hig
+ 388.400001n V_hig
+ 388.500000n V_hig
+ 388.500001n V_hig
+ 388.600000n V_hig
+ 388.600001n V_hig
+ 388.700000n V_hig
+ 388.700001n V_hig
+ 388.800000n V_hig
+ 388.800001n V_hig
+ 388.900000n V_hig
+ 388.900001n V_hig
+ 389.000000n V_hig
+ 389.000001n V_hig
+ 389.100000n V_hig
+ 389.100001n V_hig
+ 389.200000n V_hig
+ 389.200001n V_hig
+ 389.300000n V_hig
+ 389.300001n V_hig
+ 389.400000n V_hig
+ 389.400001n V_hig
+ 389.500000n V_hig
+ 389.500001n V_hig
+ 389.600000n V_hig
+ 389.600001n V_hig
+ 389.700000n V_hig
+ 389.700001n V_hig
+ 389.800000n V_hig
+ 389.800001n V_hig
+ 389.900000n V_hig
+ 389.900001n V_hig
+ 390.000000n V_hig
+ 390.000001n V_hig
+ 390.100000n V_hig
+ 390.100001n V_hig
+ 390.200000n V_hig
+ 390.200001n V_hig
+ 390.300000n V_hig
+ 390.300001n V_hig
+ 390.400000n V_hig
+ 390.400001n V_hig
+ 390.500000n V_hig
+ 390.500001n V_hig
+ 390.600000n V_hig
+ 390.600001n V_hig
+ 390.700000n V_hig
+ 390.700001n V_hig
+ 390.800000n V_hig
+ 390.800001n V_hig
+ 390.900000n V_hig
+ 390.900001n V_hig
+ 391.000000n V_hig
+ 391.000001n V_hig
+ 391.100000n V_hig
+ 391.100001n V_hig
+ 391.200000n V_hig
+ 391.200001n V_hig
+ 391.300000n V_hig
+ 391.300001n V_hig
+ 391.400000n V_hig
+ 391.400001n V_hig
+ 391.500000n V_hig
+ 391.500001n V_hig
+ 391.600000n V_hig
+ 391.600001n V_hig
+ 391.700000n V_hig
+ 391.700001n V_hig
+ 391.800000n V_hig
+ 391.800001n V_hig
+ 391.900000n V_hig
+ 391.900001n V_hig
+ 392.000000n V_hig
+ 392.000001n V_low
+ 392.100000n V_low
+ 392.100001n V_low
+ 392.200000n V_low
+ 392.200001n V_low
+ 392.300000n V_low
+ 392.300001n V_low
+ 392.400000n V_low
+ 392.400001n V_low
+ 392.500000n V_low
+ 392.500001n V_low
+ 392.600000n V_low
+ 392.600001n V_low
+ 392.700000n V_low
+ 392.700001n V_low
+ 392.800000n V_low
+ 392.800001n V_low
+ 392.900000n V_low
+ 392.900001n V_low
+ 393.000000n V_low
+ 393.000001n V_hig
+ 393.100000n V_hig
+ 393.100001n V_hig
+ 393.200000n V_hig
+ 393.200001n V_hig
+ 393.300000n V_hig
+ 393.300001n V_hig
+ 393.400000n V_hig
+ 393.400001n V_hig
+ 393.500000n V_hig
+ 393.500001n V_hig
+ 393.600000n V_hig
+ 393.600001n V_hig
+ 393.700000n V_hig
+ 393.700001n V_hig
+ 393.800000n V_hig
+ 393.800001n V_hig
+ 393.900000n V_hig
+ 393.900001n V_hig
+ 394.000000n V_hig
+ 394.000001n V_low
+ 394.100000n V_low
+ 394.100001n V_low
+ 394.200000n V_low
+ 394.200001n V_low
+ 394.300000n V_low
+ 394.300001n V_low
+ 394.400000n V_low
+ 394.400001n V_low
+ 394.500000n V_low
+ 394.500001n V_low
+ 394.600000n V_low
+ 394.600001n V_low
+ 394.700000n V_low
+ 394.700001n V_low
+ 394.800000n V_low
+ 394.800001n V_low
+ 394.900000n V_low
+ 394.900001n V_low
+ 395.000000n V_low
+ 395.000001n V_hig
+ 395.100000n V_hig
+ 395.100001n V_hig
+ 395.200000n V_hig
+ 395.200001n V_hig
+ 395.300000n V_hig
+ 395.300001n V_hig
+ 395.400000n V_hig
+ 395.400001n V_hig
+ 395.500000n V_hig
+ 395.500001n V_hig
+ 395.600000n V_hig
+ 395.600001n V_hig
+ 395.700000n V_hig
+ 395.700001n V_hig
+ 395.800000n V_hig
+ 395.800001n V_hig
+ 395.900000n V_hig
+ 395.900001n V_hig
+ 396.000000n V_hig
+ 396.000001n V_low
+ 396.100000n V_low
+ 396.100001n V_low
+ 396.200000n V_low
+ 396.200001n V_low
+ 396.300000n V_low
+ 396.300001n V_low
+ 396.400000n V_low
+ 396.400001n V_low
+ 396.500000n V_low
+ 396.500001n V_low
+ 396.600000n V_low
+ 396.600001n V_low
+ 396.700000n V_low
+ 396.700001n V_low
+ 396.800000n V_low
+ 396.800001n V_low
+ 396.900000n V_low
+ 396.900001n V_low
+ 397.000000n V_low
+ 397.000001n V_low
+ 397.100000n V_low
+ 397.100001n V_low
+ 397.200000n V_low
+ 397.200001n V_low
+ 397.300000n V_low
+ 397.300001n V_low
+ 397.400000n V_low
+ 397.400001n V_low
+ 397.500000n V_low
+ 397.500001n V_low
+ 397.600000n V_low
+ 397.600001n V_low
+ 397.700000n V_low
+ 397.700001n V_low
+ 397.800000n V_low
+ 397.800001n V_low
+ 397.900000n V_low
+ 397.900001n V_low
+ 398.000000n V_low
+ 398.000001n V_hig
+ 398.100000n V_hig
+ 398.100001n V_hig
+ 398.200000n V_hig
+ 398.200001n V_hig
+ 398.300000n V_hig
+ 398.300001n V_hig
+ 398.400000n V_hig
+ 398.400001n V_hig
+ 398.500000n V_hig
+ 398.500001n V_hig
+ 398.600000n V_hig
+ 398.600001n V_hig
+ 398.700000n V_hig
+ 398.700001n V_hig
+ 398.800000n V_hig
+ 398.800001n V_hig
+ 398.900000n V_hig
+ 398.900001n V_hig
+ 399.000000n V_hig
+ 399.000001n V_low
+ 399.100000n V_low
+ 399.100001n V_low
+ 399.200000n V_low
+ 399.200001n V_low
+ 399.300000n V_low
+ 399.300001n V_low
+ 399.400000n V_low
+ 399.400001n V_low
+ 399.500000n V_low
+ 399.500001n V_low
+ 399.600000n V_low
+ 399.600001n V_low
+ 399.700000n V_low
+ 399.700001n V_low
+ 399.800000n V_low
+ 399.800001n V_low
+ 399.900000n V_low
+ 399.900001n V_low
+ 400.000000n V_low
+ 400.000001n V_hig
+ 400.100000n V_hig
+ 400.100001n V_hig
+ 400.200000n V_hig
+ 400.200001n V_hig
+ 400.300000n V_hig
+ 400.300001n V_hig
+ 400.400000n V_hig
+ 400.400001n V_hig
+ 400.500000n V_hig
+ 400.500001n V_hig
+ 400.600000n V_hig
+ 400.600001n V_hig
+ 400.700000n V_hig
+ 400.700001n V_hig
+ 400.800000n V_hig
+ 400.800001n V_hig
+ 400.900000n V_hig
+ 400.900001n V_hig
+ 401.000000n V_hig
+ 401.000001n V_hig
+ 401.100000n V_hig
+ 401.100001n V_hig
+ 401.200000n V_hig
+ 401.200001n V_hig
+ 401.300000n V_hig
+ 401.300001n V_hig
+ 401.400000n V_hig
+ 401.400001n V_hig
+ 401.500000n V_hig
+ 401.500001n V_hig
+ 401.600000n V_hig
+ 401.600001n V_hig
+ 401.700000n V_hig
+ 401.700001n V_hig
+ 401.800000n V_hig
+ 401.800001n V_hig
+ 401.900000n V_hig
+ 401.900001n V_hig
+ 402.000000n V_hig
+ 402.000001n V_hig
+ 402.100000n V_hig
+ 402.100001n V_hig
+ 402.200000n V_hig
+ 402.200001n V_hig
+ 402.300000n V_hig
+ 402.300001n V_hig
+ 402.400000n V_hig
+ 402.400001n V_hig
+ 402.500000n V_hig
+ 402.500001n V_hig
+ 402.600000n V_hig
+ 402.600001n V_hig
+ 402.700000n V_hig
+ 402.700001n V_hig
+ 402.800000n V_hig
+ 402.800001n V_hig
+ 402.900000n V_hig
+ 402.900001n V_hig
+ 403.000000n V_hig
+ 403.000001n V_hig
+ 403.100000n V_hig
+ 403.100001n V_hig
+ 403.200000n V_hig
+ 403.200001n V_hig
+ 403.300000n V_hig
+ 403.300001n V_hig
+ 403.400000n V_hig
+ 403.400001n V_hig
+ 403.500000n V_hig
+ 403.500001n V_hig
+ 403.600000n V_hig
+ 403.600001n V_hig
+ 403.700000n V_hig
+ 403.700001n V_hig
+ 403.800000n V_hig
+ 403.800001n V_hig
+ 403.900000n V_hig
+ 403.900001n V_hig
+ 404.000000n V_hig
+ 404.000001n V_low
+ 404.100000n V_low
+ 404.100001n V_low
+ 404.200000n V_low
+ 404.200001n V_low
+ 404.300000n V_low
+ 404.300001n V_low
+ 404.400000n V_low
+ 404.400001n V_low
+ 404.500000n V_low
+ 404.500001n V_low
+ 404.600000n V_low
+ 404.600001n V_low
+ 404.700000n V_low
+ 404.700001n V_low
+ 404.800000n V_low
+ 404.800001n V_low
+ 404.900000n V_low
+ 404.900001n V_low
+ 405.000000n V_low
+ 405.000001n V_hig
+ 405.100000n V_hig
+ 405.100001n V_hig
+ 405.200000n V_hig
+ 405.200001n V_hig
+ 405.300000n V_hig
+ 405.300001n V_hig
+ 405.400000n V_hig
+ 405.400001n V_hig
+ 405.500000n V_hig
+ 405.500001n V_hig
+ 405.600000n V_hig
+ 405.600001n V_hig
+ 405.700000n V_hig
+ 405.700001n V_hig
+ 405.800000n V_hig
+ 405.800001n V_hig
+ 405.900000n V_hig
+ 405.900001n V_hig
+ 406.000000n V_hig
+ 406.000001n V_hig
+ 406.100000n V_hig
+ 406.100001n V_hig
+ 406.200000n V_hig
+ 406.200001n V_hig
+ 406.300000n V_hig
+ 406.300001n V_hig
+ 406.400000n V_hig
+ 406.400001n V_hig
+ 406.500000n V_hig
+ 406.500001n V_hig
+ 406.600000n V_hig
+ 406.600001n V_hig
+ 406.700000n V_hig
+ 406.700001n V_hig
+ 406.800000n V_hig
+ 406.800001n V_hig
+ 406.900000n V_hig
+ 406.900001n V_hig
+ 407.000000n V_hig
+ 407.000001n V_low
+ 407.100000n V_low
+ 407.100001n V_low
+ 407.200000n V_low
+ 407.200001n V_low
+ 407.300000n V_low
+ 407.300001n V_low
+ 407.400000n V_low
+ 407.400001n V_low
+ 407.500000n V_low
+ 407.500001n V_low
+ 407.600000n V_low
+ 407.600001n V_low
+ 407.700000n V_low
+ 407.700001n V_low
+ 407.800000n V_low
+ 407.800001n V_low
+ 407.900000n V_low
+ 407.900001n V_low
+ 408.000000n V_low
+ 408.000001n V_hig
+ 408.100000n V_hig
+ 408.100001n V_hig
+ 408.200000n V_hig
+ 408.200001n V_hig
+ 408.300000n V_hig
+ 408.300001n V_hig
+ 408.400000n V_hig
+ 408.400001n V_hig
+ 408.500000n V_hig
+ 408.500001n V_hig
+ 408.600000n V_hig
+ 408.600001n V_hig
+ 408.700000n V_hig
+ 408.700001n V_hig
+ 408.800000n V_hig
+ 408.800001n V_hig
+ 408.900000n V_hig
+ 408.900001n V_hig
+ 409.000000n V_hig
+ 409.000001n V_low
+ 409.100000n V_low
+ 409.100001n V_low
+ 409.200000n V_low
+ 409.200001n V_low
+ 409.300000n V_low
+ 409.300001n V_low
+ 409.400000n V_low
+ 409.400001n V_low
+ 409.500000n V_low
+ 409.500001n V_low
+ 409.600000n V_low
+ 409.600001n V_low
+ 409.700000n V_low
+ 409.700001n V_low
+ 409.800000n V_low
+ 409.800001n V_low
+ 409.900000n V_low
+ 409.900001n V_low
+ 410.000000n V_low
+ 410.000001n V_hig
+ 410.100000n V_hig
+ 410.100001n V_hig
+ 410.200000n V_hig
+ 410.200001n V_hig
+ 410.300000n V_hig
+ 410.300001n V_hig
+ 410.400000n V_hig
+ 410.400001n V_hig
+ 410.500000n V_hig
+ 410.500001n V_hig
+ 410.600000n V_hig
+ 410.600001n V_hig
+ 410.700000n V_hig
+ 410.700001n V_hig
+ 410.800000n V_hig
+ 410.800001n V_hig
+ 410.900000n V_hig
+ 410.900001n V_hig
+ 411.000000n V_hig
+ 411.000001n V_hig
+ 411.100000n V_hig
+ 411.100001n V_hig
+ 411.200000n V_hig
+ 411.200001n V_hig
+ 411.300000n V_hig
+ 411.300001n V_hig
+ 411.400000n V_hig
+ 411.400001n V_hig
+ 411.500000n V_hig
+ 411.500001n V_hig
+ 411.600000n V_hig
+ 411.600001n V_hig
+ 411.700000n V_hig
+ 411.700001n V_hig
+ 411.800000n V_hig
+ 411.800001n V_hig
+ 411.900000n V_hig
+ 411.900001n V_hig
+ 412.000000n V_hig
+ 412.000001n V_low
+ 412.100000n V_low
+ 412.100001n V_low
+ 412.200000n V_low
+ 412.200001n V_low
+ 412.300000n V_low
+ 412.300001n V_low
+ 412.400000n V_low
+ 412.400001n V_low
+ 412.500000n V_low
+ 412.500001n V_low
+ 412.600000n V_low
+ 412.600001n V_low
+ 412.700000n V_low
+ 412.700001n V_low
+ 412.800000n V_low
+ 412.800001n V_low
+ 412.900000n V_low
+ 412.900001n V_low
+ 413.000000n V_low
+ 413.000001n V_hig
+ 413.100000n V_hig
+ 413.100001n V_hig
+ 413.200000n V_hig
+ 413.200001n V_hig
+ 413.300000n V_hig
+ 413.300001n V_hig
+ 413.400000n V_hig
+ 413.400001n V_hig
+ 413.500000n V_hig
+ 413.500001n V_hig
+ 413.600000n V_hig
+ 413.600001n V_hig
+ 413.700000n V_hig
+ 413.700001n V_hig
+ 413.800000n V_hig
+ 413.800001n V_hig
+ 413.900000n V_hig
+ 413.900001n V_hig
+ 414.000000n V_hig
+ 414.000001n V_hig
+ 414.100000n V_hig
+ 414.100001n V_hig
+ 414.200000n V_hig
+ 414.200001n V_hig
+ 414.300000n V_hig
+ 414.300001n V_hig
+ 414.400000n V_hig
+ 414.400001n V_hig
+ 414.500000n V_hig
+ 414.500001n V_hig
+ 414.600000n V_hig
+ 414.600001n V_hig
+ 414.700000n V_hig
+ 414.700001n V_hig
+ 414.800000n V_hig
+ 414.800001n V_hig
+ 414.900000n V_hig
+ 414.900001n V_hig
+ 415.000000n V_hig
+ 415.000001n V_hig
+ 415.100000n V_hig
+ 415.100001n V_hig
+ 415.200000n V_hig
+ 415.200001n V_hig
+ 415.300000n V_hig
+ 415.300001n V_hig
+ 415.400000n V_hig
+ 415.400001n V_hig
+ 415.500000n V_hig
+ 415.500001n V_hig
+ 415.600000n V_hig
+ 415.600001n V_hig
+ 415.700000n V_hig
+ 415.700001n V_hig
+ 415.800000n V_hig
+ 415.800001n V_hig
+ 415.900000n V_hig
+ 415.900001n V_hig
+ 416.000000n V_hig
+ 416.000001n V_low
+ 416.100000n V_low
+ 416.100001n V_low
+ 416.200000n V_low
+ 416.200001n V_low
+ 416.300000n V_low
+ 416.300001n V_low
+ 416.400000n V_low
+ 416.400001n V_low
+ 416.500000n V_low
+ 416.500001n V_low
+ 416.600000n V_low
+ 416.600001n V_low
+ 416.700000n V_low
+ 416.700001n V_low
+ 416.800000n V_low
+ 416.800001n V_low
+ 416.900000n V_low
+ 416.900001n V_low
+ 417.000000n V_low
+ 417.000001n V_low
+ 417.100000n V_low
+ 417.100001n V_low
+ 417.200000n V_low
+ 417.200001n V_low
+ 417.300000n V_low
+ 417.300001n V_low
+ 417.400000n V_low
+ 417.400001n V_low
+ 417.500000n V_low
+ 417.500001n V_low
+ 417.600000n V_low
+ 417.600001n V_low
+ 417.700000n V_low
+ 417.700001n V_low
+ 417.800000n V_low
+ 417.800001n V_low
+ 417.900000n V_low
+ 417.900001n V_low
+ 418.000000n V_low
+ 418.000001n V_hig
+ 418.100000n V_hig
+ 418.100001n V_hig
+ 418.200000n V_hig
+ 418.200001n V_hig
+ 418.300000n V_hig
+ 418.300001n V_hig
+ 418.400000n V_hig
+ 418.400001n V_hig
+ 418.500000n V_hig
+ 418.500001n V_hig
+ 418.600000n V_hig
+ 418.600001n V_hig
+ 418.700000n V_hig
+ 418.700001n V_hig
+ 418.800000n V_hig
+ 418.800001n V_hig
+ 418.900000n V_hig
+ 418.900001n V_hig
+ 419.000000n V_hig
+ 419.000001n V_low
+ 419.100000n V_low
+ 419.100001n V_low
+ 419.200000n V_low
+ 419.200001n V_low
+ 419.300000n V_low
+ 419.300001n V_low
+ 419.400000n V_low
+ 419.400001n V_low
+ 419.500000n V_low
+ 419.500001n V_low
+ 419.600000n V_low
+ 419.600001n V_low
+ 419.700000n V_low
+ 419.700001n V_low
+ 419.800000n V_low
+ 419.800001n V_low
+ 419.900000n V_low
+ 419.900001n V_low
+ 420.000000n V_low
+ 420.000001n V_low
+ 420.100000n V_low
+ 420.100001n V_low
+ 420.200000n V_low
+ 420.200001n V_low
+ 420.300000n V_low
+ 420.300001n V_low
+ 420.400000n V_low
+ 420.400001n V_low
+ 420.500000n V_low
+ 420.500001n V_low
+ 420.600000n V_low
+ 420.600001n V_low
+ 420.700000n V_low
+ 420.700001n V_low
+ 420.800000n V_low
+ 420.800001n V_low
+ 420.900000n V_low
+ 420.900001n V_low
+ 421.000000n V_low
+ 421.000001n V_low
+ 421.100000n V_low
+ 421.100001n V_low
+ 421.200000n V_low
+ 421.200001n V_low
+ 421.300000n V_low
+ 421.300001n V_low
+ 421.400000n V_low
+ 421.400001n V_low
+ 421.500000n V_low
+ 421.500001n V_low
+ 421.600000n V_low
+ 421.600001n V_low
+ 421.700000n V_low
+ 421.700001n V_low
+ 421.800000n V_low
+ 421.800001n V_low
+ 421.900000n V_low
+ 421.900001n V_low
+ 422.000000n V_low
+ 422.000001n V_low
+ 422.100000n V_low
+ 422.100001n V_low
+ 422.200000n V_low
+ 422.200001n V_low
+ 422.300000n V_low
+ 422.300001n V_low
+ 422.400000n V_low
+ 422.400001n V_low
+ 422.500000n V_low
+ 422.500001n V_low
+ 422.600000n V_low
+ 422.600001n V_low
+ 422.700000n V_low
+ 422.700001n V_low
+ 422.800000n V_low
+ 422.800001n V_low
+ 422.900000n V_low
+ 422.900001n V_low
+ 423.000000n V_low
+ 423.000001n V_hig
+ 423.100000n V_hig
+ 423.100001n V_hig
+ 423.200000n V_hig
+ 423.200001n V_hig
+ 423.300000n V_hig
+ 423.300001n V_hig
+ 423.400000n V_hig
+ 423.400001n V_hig
+ 423.500000n V_hig
+ 423.500001n V_hig
+ 423.600000n V_hig
+ 423.600001n V_hig
+ 423.700000n V_hig
+ 423.700001n V_hig
+ 423.800000n V_hig
+ 423.800001n V_hig
+ 423.900000n V_hig
+ 423.900001n V_hig
+ 424.000000n V_hig
+ 424.000001n V_hig
+ 424.100000n V_hig
+ 424.100001n V_hig
+ 424.200000n V_hig
+ 424.200001n V_hig
+ 424.300000n V_hig
+ 424.300001n V_hig
+ 424.400000n V_hig
+ 424.400001n V_hig
+ 424.500000n V_hig
+ 424.500001n V_hig
+ 424.600000n V_hig
+ 424.600001n V_hig
+ 424.700000n V_hig
+ 424.700001n V_hig
+ 424.800000n V_hig
+ 424.800001n V_hig
+ 424.900000n V_hig
+ 424.900001n V_hig
+ 425.000000n V_hig
+ 425.000001n V_hig
+ 425.100000n V_hig
+ 425.100001n V_hig
+ 425.200000n V_hig
+ 425.200001n V_hig
+ 425.300000n V_hig
+ 425.300001n V_hig
+ 425.400000n V_hig
+ 425.400001n V_hig
+ 425.500000n V_hig
+ 425.500001n V_hig
+ 425.600000n V_hig
+ 425.600001n V_hig
+ 425.700000n V_hig
+ 425.700001n V_hig
+ 425.800000n V_hig
+ 425.800001n V_hig
+ 425.900000n V_hig
+ 425.900001n V_hig
+ 426.000000n V_hig
+ 426.000001n V_low
+ 426.100000n V_low
+ 426.100001n V_low
+ 426.200000n V_low
+ 426.200001n V_low
+ 426.300000n V_low
+ 426.300001n V_low
+ 426.400000n V_low
+ 426.400001n V_low
+ 426.500000n V_low
+ 426.500001n V_low
+ 426.600000n V_low
+ 426.600001n V_low
+ 426.700000n V_low
+ 426.700001n V_low
+ 426.800000n V_low
+ 426.800001n V_low
+ 426.900000n V_low
+ 426.900001n V_low
+ 427.000000n V_low
+ 427.000001n V_hig
+ 427.100000n V_hig
+ 427.100001n V_hig
+ 427.200000n V_hig
+ 427.200001n V_hig
+ 427.300000n V_hig
+ 427.300001n V_hig
+ 427.400000n V_hig
+ 427.400001n V_hig
+ 427.500000n V_hig
+ 427.500001n V_hig
+ 427.600000n V_hig
+ 427.600001n V_hig
+ 427.700000n V_hig
+ 427.700001n V_hig
+ 427.800000n V_hig
+ 427.800001n V_hig
+ 427.900000n V_hig
+ 427.900001n V_hig
+ 428.000000n V_hig
+ 428.000001n V_low
+ 428.100000n V_low
+ 428.100001n V_low
+ 428.200000n V_low
+ 428.200001n V_low
+ 428.300000n V_low
+ 428.300001n V_low
+ 428.400000n V_low
+ 428.400001n V_low
+ 428.500000n V_low
+ 428.500001n V_low
+ 428.600000n V_low
+ 428.600001n V_low
+ 428.700000n V_low
+ 428.700001n V_low
+ 428.800000n V_low
+ 428.800001n V_low
+ 428.900000n V_low
+ 428.900001n V_low
+ 429.000000n V_low
+ 429.000001n V_hig
+ 429.100000n V_hig
+ 429.100001n V_hig
+ 429.200000n V_hig
+ 429.200001n V_hig
+ 429.300000n V_hig
+ 429.300001n V_hig
+ 429.400000n V_hig
+ 429.400001n V_hig
+ 429.500000n V_hig
+ 429.500001n V_hig
+ 429.600000n V_hig
+ 429.600001n V_hig
+ 429.700000n V_hig
+ 429.700001n V_hig
+ 429.800000n V_hig
+ 429.800001n V_hig
+ 429.900000n V_hig
+ 429.900001n V_hig
+ 430.000000n V_hig
+ 430.000001n V_hig
+ 430.100000n V_hig
+ 430.100001n V_hig
+ 430.200000n V_hig
+ 430.200001n V_hig
+ 430.300000n V_hig
+ 430.300001n V_hig
+ 430.400000n V_hig
+ 430.400001n V_hig
+ 430.500000n V_hig
+ 430.500001n V_hig
+ 430.600000n V_hig
+ 430.600001n V_hig
+ 430.700000n V_hig
+ 430.700001n V_hig
+ 430.800000n V_hig
+ 430.800001n V_hig
+ 430.900000n V_hig
+ 430.900001n V_hig
+ 431.000000n V_hig
+ 431.000001n V_low
+ 431.100000n V_low
+ 431.100001n V_low
+ 431.200000n V_low
+ 431.200001n V_low
+ 431.300000n V_low
+ 431.300001n V_low
+ 431.400000n V_low
+ 431.400001n V_low
+ 431.500000n V_low
+ 431.500001n V_low
+ 431.600000n V_low
+ 431.600001n V_low
+ 431.700000n V_low
+ 431.700001n V_low
+ 431.800000n V_low
+ 431.800001n V_low
+ 431.900000n V_low
+ 431.900001n V_low
+ 432.000000n V_low
+ 432.000001n V_hig
+ 432.100000n V_hig
+ 432.100001n V_hig
+ 432.200000n V_hig
+ 432.200001n V_hig
+ 432.300000n V_hig
+ 432.300001n V_hig
+ 432.400000n V_hig
+ 432.400001n V_hig
+ 432.500000n V_hig
+ 432.500001n V_hig
+ 432.600000n V_hig
+ 432.600001n V_hig
+ 432.700000n V_hig
+ 432.700001n V_hig
+ 432.800000n V_hig
+ 432.800001n V_hig
+ 432.900000n V_hig
+ 432.900001n V_hig
+ 433.000000n V_hig
+ 433.000001n V_low
+ 433.100000n V_low
+ 433.100001n V_low
+ 433.200000n V_low
+ 433.200001n V_low
+ 433.300000n V_low
+ 433.300001n V_low
+ 433.400000n V_low
+ 433.400001n V_low
+ 433.500000n V_low
+ 433.500001n V_low
+ 433.600000n V_low
+ 433.600001n V_low
+ 433.700000n V_low
+ 433.700001n V_low
+ 433.800000n V_low
+ 433.800001n V_low
+ 433.900000n V_low
+ 433.900001n V_low
+ 434.000000n V_low
+ 434.000001n V_low
+ 434.100000n V_low
+ 434.100001n V_low
+ 434.200000n V_low
+ 434.200001n V_low
+ 434.300000n V_low
+ 434.300001n V_low
+ 434.400000n V_low
+ 434.400001n V_low
+ 434.500000n V_low
+ 434.500001n V_low
+ 434.600000n V_low
+ 434.600001n V_low
+ 434.700000n V_low
+ 434.700001n V_low
+ 434.800000n V_low
+ 434.800001n V_low
+ 434.900000n V_low
+ 434.900001n V_low
+ 435.000000n V_low
+ 435.000001n V_hig
+ 435.100000n V_hig
+ 435.100001n V_hig
+ 435.200000n V_hig
+ 435.200001n V_hig
+ 435.300000n V_hig
+ 435.300001n V_hig
+ 435.400000n V_hig
+ 435.400001n V_hig
+ 435.500000n V_hig
+ 435.500001n V_hig
+ 435.600000n V_hig
+ 435.600001n V_hig
+ 435.700000n V_hig
+ 435.700001n V_hig
+ 435.800000n V_hig
+ 435.800001n V_hig
+ 435.900000n V_hig
+ 435.900001n V_hig
+ 436.000000n V_hig
+ 436.000001n V_hig
+ 436.100000n V_hig
+ 436.100001n V_hig
+ 436.200000n V_hig
+ 436.200001n V_hig
+ 436.300000n V_hig
+ 436.300001n V_hig
+ 436.400000n V_hig
+ 436.400001n V_hig
+ 436.500000n V_hig
+ 436.500001n V_hig
+ 436.600000n V_hig
+ 436.600001n V_hig
+ 436.700000n V_hig
+ 436.700001n V_hig
+ 436.800000n V_hig
+ 436.800001n V_hig
+ 436.900000n V_hig
+ 436.900001n V_hig
+ 437.000000n V_hig
+ 437.000001n V_hig
+ 437.100000n V_hig
+ 437.100001n V_hig
+ 437.200000n V_hig
+ 437.200001n V_hig
+ 437.300000n V_hig
+ 437.300001n V_hig
+ 437.400000n V_hig
+ 437.400001n V_hig
+ 437.500000n V_hig
+ 437.500001n V_hig
+ 437.600000n V_hig
+ 437.600001n V_hig
+ 437.700000n V_hig
+ 437.700001n V_hig
+ 437.800000n V_hig
+ 437.800001n V_hig
+ 437.900000n V_hig
+ 437.900001n V_hig
+ 438.000000n V_hig
+ 438.000001n V_hig
+ 438.100000n V_hig
+ 438.100001n V_hig
+ 438.200000n V_hig
+ 438.200001n V_hig
+ 438.300000n V_hig
+ 438.300001n V_hig
+ 438.400000n V_hig
+ 438.400001n V_hig
+ 438.500000n V_hig
+ 438.500001n V_hig
+ 438.600000n V_hig
+ 438.600001n V_hig
+ 438.700000n V_hig
+ 438.700001n V_hig
+ 438.800000n V_hig
+ 438.800001n V_hig
+ 438.900000n V_hig
+ 438.900001n V_hig
+ 439.000000n V_hig
+ 439.000001n V_low
+ 439.100000n V_low
+ 439.100001n V_low
+ 439.200000n V_low
+ 439.200001n V_low
+ 439.300000n V_low
+ 439.300001n V_low
+ 439.400000n V_low
+ 439.400001n V_low
+ 439.500000n V_low
+ 439.500001n V_low
+ 439.600000n V_low
+ 439.600001n V_low
+ 439.700000n V_low
+ 439.700001n V_low
+ 439.800000n V_low
+ 439.800001n V_low
+ 439.900000n V_low
+ 439.900001n V_low
+ 440.000000n V_low
+ 440.000001n V_low
+ 440.100000n V_low
+ 440.100001n V_low
+ 440.200000n V_low
+ 440.200001n V_low
+ 440.300000n V_low
+ 440.300001n V_low
+ 440.400000n V_low
+ 440.400001n V_low
+ 440.500000n V_low
+ 440.500001n V_low
+ 440.600000n V_low
+ 440.600001n V_low
+ 440.700000n V_low
+ 440.700001n V_low
+ 440.800000n V_low
+ 440.800001n V_low
+ 440.900000n V_low
+ 440.900001n V_low
+ 441.000000n V_low
+ 441.000001n V_low
+ 441.100000n V_low
+ 441.100001n V_low
+ 441.200000n V_low
+ 441.200001n V_low
+ 441.300000n V_low
+ 441.300001n V_low
+ 441.400000n V_low
+ 441.400001n V_low
+ 441.500000n V_low
+ 441.500001n V_low
+ 441.600000n V_low
+ 441.600001n V_low
+ 441.700000n V_low
+ 441.700001n V_low
+ 441.800000n V_low
+ 441.800001n V_low
+ 441.900000n V_low
+ 441.900001n V_low
+ 442.000000n V_low
+ 442.000001n V_hig
+ 442.100000n V_hig
+ 442.100001n V_hig
+ 442.200000n V_hig
+ 442.200001n V_hig
+ 442.300000n V_hig
+ 442.300001n V_hig
+ 442.400000n V_hig
+ 442.400001n V_hig
+ 442.500000n V_hig
+ 442.500001n V_hig
+ 442.600000n V_hig
+ 442.600001n V_hig
+ 442.700000n V_hig
+ 442.700001n V_hig
+ 442.800000n V_hig
+ 442.800001n V_hig
+ 442.900000n V_hig
+ 442.900001n V_hig
+ 443.000000n V_hig
+ 443.000001n V_low
+ 443.100000n V_low
+ 443.100001n V_low
+ 443.200000n V_low
+ 443.200001n V_low
+ 443.300000n V_low
+ 443.300001n V_low
+ 443.400000n V_low
+ 443.400001n V_low
+ 443.500000n V_low
+ 443.500001n V_low
+ 443.600000n V_low
+ 443.600001n V_low
+ 443.700000n V_low
+ 443.700001n V_low
+ 443.800000n V_low
+ 443.800001n V_low
+ 443.900000n V_low
+ 443.900001n V_low
+ 444.000000n V_low
+ 444.000001n V_hig
+ 444.100000n V_hig
+ 444.100001n V_hig
+ 444.200000n V_hig
+ 444.200001n V_hig
+ 444.300000n V_hig
+ 444.300001n V_hig
+ 444.400000n V_hig
+ 444.400001n V_hig
+ 444.500000n V_hig
+ 444.500001n V_hig
+ 444.600000n V_hig
+ 444.600001n V_hig
+ 444.700000n V_hig
+ 444.700001n V_hig
+ 444.800000n V_hig
+ 444.800001n V_hig
+ 444.900000n V_hig
+ 444.900001n V_hig
+ 445.000000n V_hig
+ 445.000001n V_hig
+ 445.100000n V_hig
+ 445.100001n V_hig
+ 445.200000n V_hig
+ 445.200001n V_hig
+ 445.300000n V_hig
+ 445.300001n V_hig
+ 445.400000n V_hig
+ 445.400001n V_hig
+ 445.500000n V_hig
+ 445.500001n V_hig
+ 445.600000n V_hig
+ 445.600001n V_hig
+ 445.700000n V_hig
+ 445.700001n V_hig
+ 445.800000n V_hig
+ 445.800001n V_hig
+ 445.900000n V_hig
+ 445.900001n V_hig
+ 446.000000n V_hig
+ 446.000001n V_low
+ 446.100000n V_low
+ 446.100001n V_low
+ 446.200000n V_low
+ 446.200001n V_low
+ 446.300000n V_low
+ 446.300001n V_low
+ 446.400000n V_low
+ 446.400001n V_low
+ 446.500000n V_low
+ 446.500001n V_low
+ 446.600000n V_low
+ 446.600001n V_low
+ 446.700000n V_low
+ 446.700001n V_low
+ 446.800000n V_low
+ 446.800001n V_low
+ 446.900000n V_low
+ 446.900001n V_low
+ 447.000000n V_low
+ 447.000001n V_low
+ 447.100000n V_low
+ 447.100001n V_low
+ 447.200000n V_low
+ 447.200001n V_low
+ 447.300000n V_low
+ 447.300001n V_low
+ 447.400000n V_low
+ 447.400001n V_low
+ 447.500000n V_low
+ 447.500001n V_low
+ 447.600000n V_low
+ 447.600001n V_low
+ 447.700000n V_low
+ 447.700001n V_low
+ 447.800000n V_low
+ 447.800001n V_low
+ 447.900000n V_low
+ 447.900001n V_low
+ 448.000000n V_low
+ 448.000001n V_low
+ 448.100000n V_low
+ 448.100001n V_low
+ 448.200000n V_low
+ 448.200001n V_low
+ 448.300000n V_low
+ 448.300001n V_low
+ 448.400000n V_low
+ 448.400001n V_low
+ 448.500000n V_low
+ 448.500001n V_low
+ 448.600000n V_low
+ 448.600001n V_low
+ 448.700000n V_low
+ 448.700001n V_low
+ 448.800000n V_low
+ 448.800001n V_low
+ 448.900000n V_low
+ 448.900001n V_low
+ 449.000000n V_low
+ 449.000001n V_low
+ 449.100000n V_low
+ 449.100001n V_low
+ 449.200000n V_low
+ 449.200001n V_low
+ 449.300000n V_low
+ 449.300001n V_low
+ 449.400000n V_low
+ 449.400001n V_low
+ 449.500000n V_low
+ 449.500001n V_low
+ 449.600000n V_low
+ 449.600001n V_low
+ 449.700000n V_low
+ 449.700001n V_low
+ 449.800000n V_low
+ 449.800001n V_low
+ 449.900000n V_low
+ 449.900001n V_low
+ 450.000000n V_low
+ 450.000001n V_low
+ 450.100000n V_low
+ 450.100001n V_low
+ 450.200000n V_low
+ 450.200001n V_low
+ 450.300000n V_low
+ 450.300001n V_low
+ 450.400000n V_low
+ 450.400001n V_low
+ 450.500000n V_low
+ 450.500001n V_low
+ 450.600000n V_low
+ 450.600001n V_low
+ 450.700000n V_low
+ 450.700001n V_low
+ 450.800000n V_low
+ 450.800001n V_low
+ 450.900000n V_low
+ 450.900001n V_low
+ 451.000000n V_low
+ 451.000001n V_hig
+ 451.100000n V_hig
+ 451.100001n V_hig
+ 451.200000n V_hig
+ 451.200001n V_hig
+ 451.300000n V_hig
+ 451.300001n V_hig
+ 451.400000n V_hig
+ 451.400001n V_hig
+ 451.500000n V_hig
+ 451.500001n V_hig
+ 451.600000n V_hig
+ 451.600001n V_hig
+ 451.700000n V_hig
+ 451.700001n V_hig
+ 451.800000n V_hig
+ 451.800001n V_hig
+ 451.900000n V_hig
+ 451.900001n V_hig
+ 452.000000n V_hig
+ 452.000001n V_hig
+ 452.100000n V_hig
+ 452.100001n V_hig
+ 452.200000n V_hig
+ 452.200001n V_hig
+ 452.300000n V_hig
+ 452.300001n V_hig
+ 452.400000n V_hig
+ 452.400001n V_hig
+ 452.500000n V_hig
+ 452.500001n V_hig
+ 452.600000n V_hig
+ 452.600001n V_hig
+ 452.700000n V_hig
+ 452.700001n V_hig
+ 452.800000n V_hig
+ 452.800001n V_hig
+ 452.900000n V_hig
+ 452.900001n V_hig
+ 453.000000n V_hig
+ 453.000001n V_low
+ 453.100000n V_low
+ 453.100001n V_low
+ 453.200000n V_low
+ 453.200001n V_low
+ 453.300000n V_low
+ 453.300001n V_low
+ 453.400000n V_low
+ 453.400001n V_low
+ 453.500000n V_low
+ 453.500001n V_low
+ 453.600000n V_low
+ 453.600001n V_low
+ 453.700000n V_low
+ 453.700001n V_low
+ 453.800000n V_low
+ 453.800001n V_low
+ 453.900000n V_low
+ 453.900001n V_low
+ 454.000000n V_low
+ 454.000001n V_low
+ 454.100000n V_low
+ 454.100001n V_low
+ 454.200000n V_low
+ 454.200001n V_low
+ 454.300000n V_low
+ 454.300001n V_low
+ 454.400000n V_low
+ 454.400001n V_low
+ 454.500000n V_low
+ 454.500001n V_low
+ 454.600000n V_low
+ 454.600001n V_low
+ 454.700000n V_low
+ 454.700001n V_low
+ 454.800000n V_low
+ 454.800001n V_low
+ 454.900000n V_low
+ 454.900001n V_low
+ 455.000000n V_low
+ 455.000001n V_low
+ 455.100000n V_low
+ 455.100001n V_low
+ 455.200000n V_low
+ 455.200001n V_low
+ 455.300000n V_low
+ 455.300001n V_low
+ 455.400000n V_low
+ 455.400001n V_low
+ 455.500000n V_low
+ 455.500001n V_low
+ 455.600000n V_low
+ 455.600001n V_low
+ 455.700000n V_low
+ 455.700001n V_low
+ 455.800000n V_low
+ 455.800001n V_low
+ 455.900000n V_low
+ 455.900001n V_low
+ 456.000000n V_low
+ 456.000001n V_low
+ 456.100000n V_low
+ 456.100001n V_low
+ 456.200000n V_low
+ 456.200001n V_low
+ 456.300000n V_low
+ 456.300001n V_low
+ 456.400000n V_low
+ 456.400001n V_low
+ 456.500000n V_low
+ 456.500001n V_low
+ 456.600000n V_low
+ 456.600001n V_low
+ 456.700000n V_low
+ 456.700001n V_low
+ 456.800000n V_low
+ 456.800001n V_low
+ 456.900000n V_low
+ 456.900001n V_low
+ 457.000000n V_low
+ 457.000001n V_hig
+ 457.100000n V_hig
+ 457.100001n V_hig
+ 457.200000n V_hig
+ 457.200001n V_hig
+ 457.300000n V_hig
+ 457.300001n V_hig
+ 457.400000n V_hig
+ 457.400001n V_hig
+ 457.500000n V_hig
+ 457.500001n V_hig
+ 457.600000n V_hig
+ 457.600001n V_hig
+ 457.700000n V_hig
+ 457.700001n V_hig
+ 457.800000n V_hig
+ 457.800001n V_hig
+ 457.900000n V_hig
+ 457.900001n V_hig
+ 458.000000n V_hig
+ 458.000001n V_low
+ 458.100000n V_low
+ 458.100001n V_low
+ 458.200000n V_low
+ 458.200001n V_low
+ 458.300000n V_low
+ 458.300001n V_low
+ 458.400000n V_low
+ 458.400001n V_low
+ 458.500000n V_low
+ 458.500001n V_low
+ 458.600000n V_low
+ 458.600001n V_low
+ 458.700000n V_low
+ 458.700001n V_low
+ 458.800000n V_low
+ 458.800001n V_low
+ 458.900000n V_low
+ 458.900001n V_low
+ 459.000000n V_low
+ 459.000001n V_hig
+ 459.100000n V_hig
+ 459.100001n V_hig
+ 459.200000n V_hig
+ 459.200001n V_hig
+ 459.300000n V_hig
+ 459.300001n V_hig
+ 459.400000n V_hig
+ 459.400001n V_hig
+ 459.500000n V_hig
+ 459.500001n V_hig
+ 459.600000n V_hig
+ 459.600001n V_hig
+ 459.700000n V_hig
+ 459.700001n V_hig
+ 459.800000n V_hig
+ 459.800001n V_hig
+ 459.900000n V_hig
+ 459.900001n V_hig
+ 460.000000n V_hig
+ 460.000001n V_low
+ 460.100000n V_low
+ 460.100001n V_low
+ 460.200000n V_low
+ 460.200001n V_low
+ 460.300000n V_low
+ 460.300001n V_low
+ 460.400000n V_low
+ 460.400001n V_low
+ 460.500000n V_low
+ 460.500001n V_low
+ 460.600000n V_low
+ 460.600001n V_low
+ 460.700000n V_low
+ 460.700001n V_low
+ 460.800000n V_low
+ 460.800001n V_low
+ 460.900000n V_low
+ 460.900001n V_low
+ 461.000000n V_low
+ 461.000001n V_low
+ 461.100000n V_low
+ 461.100001n V_low
+ 461.200000n V_low
+ 461.200001n V_low
+ 461.300000n V_low
+ 461.300001n V_low
+ 461.400000n V_low
+ 461.400001n V_low
+ 461.500000n V_low
+ 461.500001n V_low
+ 461.600000n V_low
+ 461.600001n V_low
+ 461.700000n V_low
+ 461.700001n V_low
+ 461.800000n V_low
+ 461.800001n V_low
+ 461.900000n V_low
+ 461.900001n V_low
+ 462.000000n V_low
+ 462.000001n V_hig
+ 462.100000n V_hig
+ 462.100001n V_hig
+ 462.200000n V_hig
+ 462.200001n V_hig
+ 462.300000n V_hig
+ 462.300001n V_hig
+ 462.400000n V_hig
+ 462.400001n V_hig
+ 462.500000n V_hig
+ 462.500001n V_hig
+ 462.600000n V_hig
+ 462.600001n V_hig
+ 462.700000n V_hig
+ 462.700001n V_hig
+ 462.800000n V_hig
+ 462.800001n V_hig
+ 462.900000n V_hig
+ 462.900001n V_hig
+ 463.000000n V_hig
+ 463.000001n V_low
+ 463.100000n V_low
+ 463.100001n V_low
+ 463.200000n V_low
+ 463.200001n V_low
+ 463.300000n V_low
+ 463.300001n V_low
+ 463.400000n V_low
+ 463.400001n V_low
+ 463.500000n V_low
+ 463.500001n V_low
+ 463.600000n V_low
+ 463.600001n V_low
+ 463.700000n V_low
+ 463.700001n V_low
+ 463.800000n V_low
+ 463.800001n V_low
+ 463.900000n V_low
+ 463.900001n V_low
+ 464.000000n V_low
+ 464.000001n V_low
+ 464.100000n V_low
+ 464.100001n V_low
+ 464.200000n V_low
+ 464.200001n V_low
+ 464.300000n V_low
+ 464.300001n V_low
+ 464.400000n V_low
+ 464.400001n V_low
+ 464.500000n V_low
+ 464.500001n V_low
+ 464.600000n V_low
+ 464.600001n V_low
+ 464.700000n V_low
+ 464.700001n V_low
+ 464.800000n V_low
+ 464.800001n V_low
+ 464.900000n V_low
+ 464.900001n V_low
+ 465.000000n V_low
+ 465.000001n V_hig
+ 465.100000n V_hig
+ 465.100001n V_hig
+ 465.200000n V_hig
+ 465.200001n V_hig
+ 465.300000n V_hig
+ 465.300001n V_hig
+ 465.400000n V_hig
+ 465.400001n V_hig
+ 465.500000n V_hig
+ 465.500001n V_hig
+ 465.600000n V_hig
+ 465.600001n V_hig
+ 465.700000n V_hig
+ 465.700001n V_hig
+ 465.800000n V_hig
+ 465.800001n V_hig
+ 465.900000n V_hig
+ 465.900001n V_hig
+ 466.000000n V_hig
+ 466.000001n V_low
+ 466.100000n V_low
+ 466.100001n V_low
+ 466.200000n V_low
+ 466.200001n V_low
+ 466.300000n V_low
+ 466.300001n V_low
+ 466.400000n V_low
+ 466.400001n V_low
+ 466.500000n V_low
+ 466.500001n V_low
+ 466.600000n V_low
+ 466.600001n V_low
+ 466.700000n V_low
+ 466.700001n V_low
+ 466.800000n V_low
+ 466.800001n V_low
+ 466.900000n V_low
+ 466.900001n V_low
+ 467.000000n V_low
+ 467.000001n V_hig
+ 467.100000n V_hig
+ 467.100001n V_hig
+ 467.200000n V_hig
+ 467.200001n V_hig
+ 467.300000n V_hig
+ 467.300001n V_hig
+ 467.400000n V_hig
+ 467.400001n V_hig
+ 467.500000n V_hig
+ 467.500001n V_hig
+ 467.600000n V_hig
+ 467.600001n V_hig
+ 467.700000n V_hig
+ 467.700001n V_hig
+ 467.800000n V_hig
+ 467.800001n V_hig
+ 467.900000n V_hig
+ 467.900001n V_hig
+ 468.000000n V_hig
+ 468.000001n V_low
+ 468.100000n V_low
+ 468.100001n V_low
+ 468.200000n V_low
+ 468.200001n V_low
+ 468.300000n V_low
+ 468.300001n V_low
+ 468.400000n V_low
+ 468.400001n V_low
+ 468.500000n V_low
+ 468.500001n V_low
+ 468.600000n V_low
+ 468.600001n V_low
+ 468.700000n V_low
+ 468.700001n V_low
+ 468.800000n V_low
+ 468.800001n V_low
+ 468.900000n V_low
+ 468.900001n V_low
+ 469.000000n V_low
+ 469.000001n V_low
+ 469.100000n V_low
+ 469.100001n V_low
+ 469.200000n V_low
+ 469.200001n V_low
+ 469.300000n V_low
+ 469.300001n V_low
+ 469.400000n V_low
+ 469.400001n V_low
+ 469.500000n V_low
+ 469.500001n V_low
+ 469.600000n V_low
+ 469.600001n V_low
+ 469.700000n V_low
+ 469.700001n V_low
+ 469.800000n V_low
+ 469.800001n V_low
+ 469.900000n V_low
+ 469.900001n V_low
+ 470.000000n V_low
+ 470.000001n V_low
+ 470.100000n V_low
+ 470.100001n V_low
+ 470.200000n V_low
+ 470.200001n V_low
+ 470.300000n V_low
+ 470.300001n V_low
+ 470.400000n V_low
+ 470.400001n V_low
+ 470.500000n V_low
+ 470.500001n V_low
+ 470.600000n V_low
+ 470.600001n V_low
+ 470.700000n V_low
+ 470.700001n V_low
+ 470.800000n V_low
+ 470.800001n V_low
+ 470.900000n V_low
+ 470.900001n V_low
+ 471.000000n V_low
+ 471.000001n V_hig
+ 471.100000n V_hig
+ 471.100001n V_hig
+ 471.200000n V_hig
+ 471.200001n V_hig
+ 471.300000n V_hig
+ 471.300001n V_hig
+ 471.400000n V_hig
+ 471.400001n V_hig
+ 471.500000n V_hig
+ 471.500001n V_hig
+ 471.600000n V_hig
+ 471.600001n V_hig
+ 471.700000n V_hig
+ 471.700001n V_hig
+ 471.800000n V_hig
+ 471.800001n V_hig
+ 471.900000n V_hig
+ 471.900001n V_hig
+ 472.000000n V_hig
+ 472.000001n V_hig
+ 472.100000n V_hig
+ 472.100001n V_hig
+ 472.200000n V_hig
+ 472.200001n V_hig
+ 472.300000n V_hig
+ 472.300001n V_hig
+ 472.400000n V_hig
+ 472.400001n V_hig
+ 472.500000n V_hig
+ 472.500001n V_hig
+ 472.600000n V_hig
+ 472.600001n V_hig
+ 472.700000n V_hig
+ 472.700001n V_hig
+ 472.800000n V_hig
+ 472.800001n V_hig
+ 472.900000n V_hig
+ 472.900001n V_hig
+ 473.000000n V_hig
+ 473.000001n V_low
+ 473.100000n V_low
+ 473.100001n V_low
+ 473.200000n V_low
+ 473.200001n V_low
+ 473.300000n V_low
+ 473.300001n V_low
+ 473.400000n V_low
+ 473.400001n V_low
+ 473.500000n V_low
+ 473.500001n V_low
+ 473.600000n V_low
+ 473.600001n V_low
+ 473.700000n V_low
+ 473.700001n V_low
+ 473.800000n V_low
+ 473.800001n V_low
+ 473.900000n V_low
+ 473.900001n V_low
+ 474.000000n V_low
+ 474.000001n V_hig
+ 474.100000n V_hig
+ 474.100001n V_hig
+ 474.200000n V_hig
+ 474.200001n V_hig
+ 474.300000n V_hig
+ 474.300001n V_hig
+ 474.400000n V_hig
+ 474.400001n V_hig
+ 474.500000n V_hig
+ 474.500001n V_hig
+ 474.600000n V_hig
+ 474.600001n V_hig
+ 474.700000n V_hig
+ 474.700001n V_hig
+ 474.800000n V_hig
+ 474.800001n V_hig
+ 474.900000n V_hig
+ 474.900001n V_hig
+ 475.000000n V_hig
+ 475.000001n V_hig
+ 475.100000n V_hig
+ 475.100001n V_hig
+ 475.200000n V_hig
+ 475.200001n V_hig
+ 475.300000n V_hig
+ 475.300001n V_hig
+ 475.400000n V_hig
+ 475.400001n V_hig
+ 475.500000n V_hig
+ 475.500001n V_hig
+ 475.600000n V_hig
+ 475.600001n V_hig
+ 475.700000n V_hig
+ 475.700001n V_hig
+ 475.800000n V_hig
+ 475.800001n V_hig
+ 475.900000n V_hig
+ 475.900001n V_hig
+ 476.000000n V_hig
+ 476.000001n V_hig
+ 476.100000n V_hig
+ 476.100001n V_hig
+ 476.200000n V_hig
+ 476.200001n V_hig
+ 476.300000n V_hig
+ 476.300001n V_hig
+ 476.400000n V_hig
+ 476.400001n V_hig
+ 476.500000n V_hig
+ 476.500001n V_hig
+ 476.600000n V_hig
+ 476.600001n V_hig
+ 476.700000n V_hig
+ 476.700001n V_hig
+ 476.800000n V_hig
+ 476.800001n V_hig
+ 476.900000n V_hig
+ 476.900001n V_hig
+ 477.000000n V_hig
+ 477.000001n V_low
+ 477.100000n V_low
+ 477.100001n V_low
+ 477.200000n V_low
+ 477.200001n V_low
+ 477.300000n V_low
+ 477.300001n V_low
+ 477.400000n V_low
+ 477.400001n V_low
+ 477.500000n V_low
+ 477.500001n V_low
+ 477.600000n V_low
+ 477.600001n V_low
+ 477.700000n V_low
+ 477.700001n V_low
+ 477.800000n V_low
+ 477.800001n V_low
+ 477.900000n V_low
+ 477.900001n V_low
+ 478.000000n V_low
+ 478.000001n V_hig
+ 478.100000n V_hig
+ 478.100001n V_hig
+ 478.200000n V_hig
+ 478.200001n V_hig
+ 478.300000n V_hig
+ 478.300001n V_hig
+ 478.400000n V_hig
+ 478.400001n V_hig
+ 478.500000n V_hig
+ 478.500001n V_hig
+ 478.600000n V_hig
+ 478.600001n V_hig
+ 478.700000n V_hig
+ 478.700001n V_hig
+ 478.800000n V_hig
+ 478.800001n V_hig
+ 478.900000n V_hig
+ 478.900001n V_hig
+ 479.000000n V_hig
+ 479.000001n V_low
+ 479.100000n V_low
+ 479.100001n V_low
+ 479.200000n V_low
+ 479.200001n V_low
+ 479.300000n V_low
+ 479.300001n V_low
+ 479.400000n V_low
+ 479.400001n V_low
+ 479.500000n V_low
+ 479.500001n V_low
+ 479.600000n V_low
+ 479.600001n V_low
+ 479.700000n V_low
+ 479.700001n V_low
+ 479.800000n V_low
+ 479.800001n V_low
+ 479.900000n V_low
+ 479.900001n V_low
+ 480.000000n V_low
+ 480.000001n V_low
+ 480.100000n V_low
+ 480.100001n V_low
+ 480.200000n V_low
+ 480.200001n V_low
+ 480.300000n V_low
+ 480.300001n V_low
+ 480.400000n V_low
+ 480.400001n V_low
+ 480.500000n V_low
+ 480.500001n V_low
+ 480.600000n V_low
+ 480.600001n V_low
+ 480.700000n V_low
+ 480.700001n V_low
+ 480.800000n V_low
+ 480.800001n V_low
+ 480.900000n V_low
+ 480.900001n V_low
+ 481.000000n V_low
+ 481.000001n V_low
+ 481.100000n V_low
+ 481.100001n V_low
+ 481.200000n V_low
+ 481.200001n V_low
+ 481.300000n V_low
+ 481.300001n V_low
+ 481.400000n V_low
+ 481.400001n V_low
+ 481.500000n V_low
+ 481.500001n V_low
+ 481.600000n V_low
+ 481.600001n V_low
+ 481.700000n V_low
+ 481.700001n V_low
+ 481.800000n V_low
+ 481.800001n V_low
+ 481.900000n V_low
+ 481.900001n V_low
+ 482.000000n V_low
+ 482.000001n V_low
+ 482.100000n V_low
+ 482.100001n V_low
+ 482.200000n V_low
+ 482.200001n V_low
+ 482.300000n V_low
+ 482.300001n V_low
+ 482.400000n V_low
+ 482.400001n V_low
+ 482.500000n V_low
+ 482.500001n V_low
+ 482.600000n V_low
+ 482.600001n V_low
+ 482.700000n V_low
+ 482.700001n V_low
+ 482.800000n V_low
+ 482.800001n V_low
+ 482.900000n V_low
+ 482.900001n V_low
+ 483.000000n V_low
+ 483.000001n V_low
+ 483.100000n V_low
+ 483.100001n V_low
+ 483.200000n V_low
+ 483.200001n V_low
+ 483.300000n V_low
+ 483.300001n V_low
+ 483.400000n V_low
+ 483.400001n V_low
+ 483.500000n V_low
+ 483.500001n V_low
+ 483.600000n V_low
+ 483.600001n V_low
+ 483.700000n V_low
+ 483.700001n V_low
+ 483.800000n V_low
+ 483.800001n V_low
+ 483.900000n V_low
+ 483.900001n V_low
+ 484.000000n V_low
+ 484.000001n V_hig
+ 484.100000n V_hig
+ 484.100001n V_hig
+ 484.200000n V_hig
+ 484.200001n V_hig
+ 484.300000n V_hig
+ 484.300001n V_hig
+ 484.400000n V_hig
+ 484.400001n V_hig
+ 484.500000n V_hig
+ 484.500001n V_hig
+ 484.600000n V_hig
+ 484.600001n V_hig
+ 484.700000n V_hig
+ 484.700001n V_hig
+ 484.800000n V_hig
+ 484.800001n V_hig
+ 484.900000n V_hig
+ 484.900001n V_hig
+ 485.000000n V_hig
+ 485.000001n V_low
+ 485.100000n V_low
+ 485.100001n V_low
+ 485.200000n V_low
+ 485.200001n V_low
+ 485.300000n V_low
+ 485.300001n V_low
+ 485.400000n V_low
+ 485.400001n V_low
+ 485.500000n V_low
+ 485.500001n V_low
+ 485.600000n V_low
+ 485.600001n V_low
+ 485.700000n V_low
+ 485.700001n V_low
+ 485.800000n V_low
+ 485.800001n V_low
+ 485.900000n V_low
+ 485.900001n V_low
+ 486.000000n V_low
+ 486.000001n V_hig
+ 486.100000n V_hig
+ 486.100001n V_hig
+ 486.200000n V_hig
+ 486.200001n V_hig
+ 486.300000n V_hig
+ 486.300001n V_hig
+ 486.400000n V_hig
+ 486.400001n V_hig
+ 486.500000n V_hig
+ 486.500001n V_hig
+ 486.600000n V_hig
+ 486.600001n V_hig
+ 486.700000n V_hig
+ 486.700001n V_hig
+ 486.800000n V_hig
+ 486.800001n V_hig
+ 486.900000n V_hig
+ 486.900001n V_hig
+ 487.000000n V_hig
+ 487.000001n V_hig
+ 487.100000n V_hig
+ 487.100001n V_hig
+ 487.200000n V_hig
+ 487.200001n V_hig
+ 487.300000n V_hig
+ 487.300001n V_hig
+ 487.400000n V_hig
+ 487.400001n V_hig
+ 487.500000n V_hig
+ 487.500001n V_hig
+ 487.600000n V_hig
+ 487.600001n V_hig
+ 487.700000n V_hig
+ 487.700001n V_hig
+ 487.800000n V_hig
+ 487.800001n V_hig
+ 487.900000n V_hig
+ 487.900001n V_hig
+ 488.000000n V_hig
+ 488.000001n V_low
+ 488.100000n V_low
+ 488.100001n V_low
+ 488.200000n V_low
+ 488.200001n V_low
+ 488.300000n V_low
+ 488.300001n V_low
+ 488.400000n V_low
+ 488.400001n V_low
+ 488.500000n V_low
+ 488.500001n V_low
+ 488.600000n V_low
+ 488.600001n V_low
+ 488.700000n V_low
+ 488.700001n V_low
+ 488.800000n V_low
+ 488.800001n V_low
+ 488.900000n V_low
+ 488.900001n V_low
+ 489.000000n V_low
+ 489.000001n V_low
+ 489.100000n V_low
+ 489.100001n V_low
+ 489.200000n V_low
+ 489.200001n V_low
+ 489.300000n V_low
+ 489.300001n V_low
+ 489.400000n V_low
+ 489.400001n V_low
+ 489.500000n V_low
+ 489.500001n V_low
+ 489.600000n V_low
+ 489.600001n V_low
+ 489.700000n V_low
+ 489.700001n V_low
+ 489.800000n V_low
+ 489.800001n V_low
+ 489.900000n V_low
+ 489.900001n V_low
+ 490.000000n V_low
+ 490.000001n V_hig
+ 490.100000n V_hig
+ 490.100001n V_hig
+ 490.200000n V_hig
+ 490.200001n V_hig
+ 490.300000n V_hig
+ 490.300001n V_hig
+ 490.400000n V_hig
+ 490.400001n V_hig
+ 490.500000n V_hig
+ 490.500001n V_hig
+ 490.600000n V_hig
+ 490.600001n V_hig
+ 490.700000n V_hig
+ 490.700001n V_hig
+ 490.800000n V_hig
+ 490.800001n V_hig
+ 490.900000n V_hig
+ 490.900001n V_hig
+ 491.000000n V_hig
+ 491.000001n V_hig
+ 491.100000n V_hig
+ 491.100001n V_hig
+ 491.200000n V_hig
+ 491.200001n V_hig
+ 491.300000n V_hig
+ 491.300001n V_hig
+ 491.400000n V_hig
+ 491.400001n V_hig
+ 491.500000n V_hig
+ 491.500001n V_hig
+ 491.600000n V_hig
+ 491.600001n V_hig
+ 491.700000n V_hig
+ 491.700001n V_hig
+ 491.800000n V_hig
+ 491.800001n V_hig
+ 491.900000n V_hig
+ 491.900001n V_hig
+ 492.000000n V_hig
+ 492.000001n V_hig
+ 492.100000n V_hig
+ 492.100001n V_hig
+ 492.200000n V_hig
+ 492.200001n V_hig
+ 492.300000n V_hig
+ 492.300001n V_hig
+ 492.400000n V_hig
+ 492.400001n V_hig
+ 492.500000n V_hig
+ 492.500001n V_hig
+ 492.600000n V_hig
+ 492.600001n V_hig
+ 492.700000n V_hig
+ 492.700001n V_hig
+ 492.800000n V_hig
+ 492.800001n V_hig
+ 492.900000n V_hig
+ 492.900001n V_hig
+ 493.000000n V_hig
+ 493.000001n V_low
+ 493.100000n V_low
+ 493.100001n V_low
+ 493.200000n V_low
+ 493.200001n V_low
+ 493.300000n V_low
+ 493.300001n V_low
+ 493.400000n V_low
+ 493.400001n V_low
+ 493.500000n V_low
+ 493.500001n V_low
+ 493.600000n V_low
+ 493.600001n V_low
+ 493.700000n V_low
+ 493.700001n V_low
+ 493.800000n V_low
+ 493.800001n V_low
+ 493.900000n V_low
+ 493.900001n V_low
+ 494.000000n V_low
+ 494.000001n V_low
+ 494.100000n V_low
+ 494.100001n V_low
+ 494.200000n V_low
+ 494.200001n V_low
+ 494.300000n V_low
+ 494.300001n V_low
+ 494.400000n V_low
+ 494.400001n V_low
+ 494.500000n V_low
+ 494.500001n V_low
+ 494.600000n V_low
+ 494.600001n V_low
+ 494.700000n V_low
+ 494.700001n V_low
+ 494.800000n V_low
+ 494.800001n V_low
+ 494.900000n V_low
+ 494.900001n V_low
+ 495.000000n V_low
+ 495.000001n V_low
+ 495.100000n V_low
+ 495.100001n V_low
+ 495.200000n V_low
+ 495.200001n V_low
+ 495.300000n V_low
+ 495.300001n V_low
+ 495.400000n V_low
+ 495.400001n V_low
+ 495.500000n V_low
+ 495.500001n V_low
+ 495.600000n V_low
+ 495.600001n V_low
+ 495.700000n V_low
+ 495.700001n V_low
+ 495.800000n V_low
+ 495.800001n V_low
+ 495.900000n V_low
+ 495.900001n V_low
+ 496.000000n V_low
+ 496.000001n V_hig
+ 496.100000n V_hig
+ 496.100001n V_hig
+ 496.200000n V_hig
+ 496.200001n V_hig
+ 496.300000n V_hig
+ 496.300001n V_hig
+ 496.400000n V_hig
+ 496.400001n V_hig
+ 496.500000n V_hig
+ 496.500001n V_hig
+ 496.600000n V_hig
+ 496.600001n V_hig
+ 496.700000n V_hig
+ 496.700001n V_hig
+ 496.800000n V_hig
+ 496.800001n V_hig
+ 496.900000n V_hig
+ 496.900001n V_hig
+ 497.000000n V_hig
+ 497.000001n V_hig
+ 497.100000n V_hig
+ 497.100001n V_hig
+ 497.200000n V_hig
+ 497.200001n V_hig
+ 497.300000n V_hig
+ 497.300001n V_hig
+ 497.400000n V_hig
+ 497.400001n V_hig
+ 497.500000n V_hig
+ 497.500001n V_hig
+ 497.600000n V_hig
+ 497.600001n V_hig
+ 497.700000n V_hig
+ 497.700001n V_hig
+ 497.800000n V_hig
+ 497.800001n V_hig
+ 497.900000n V_hig
+ 497.900001n V_hig
+ 498.000000n V_hig
+ 498.000001n V_low
+ 498.100000n V_low
+ 498.100001n V_low
+ 498.200000n V_low
+ 498.200001n V_low
+ 498.300000n V_low
+ 498.300001n V_low
+ 498.400000n V_low
+ 498.400001n V_low
+ 498.500000n V_low
+ 498.500001n V_low
+ 498.600000n V_low
+ 498.600001n V_low
+ 498.700000n V_low
+ 498.700001n V_low
+ 498.800000n V_low
+ 498.800001n V_low
+ 498.900000n V_low
+ 498.900001n V_low
+ 499.000000n V_low
+ 499.000001n V_low
+ 499.100000n V_low
+ 499.100001n V_low
+ 499.200000n V_low
+ 499.200001n V_low
+ 499.300000n V_low
+ 499.300001n V_low
+ 499.400000n V_low
+ 499.400001n V_low
+ 499.500000n V_low
+ 499.500001n V_low
+ 499.600000n V_low
+ 499.600001n V_low
+ 499.700000n V_low
+ 499.700001n V_low
+ 499.800000n V_low
+ 499.800001n V_low
+ 499.900000n V_low
+ 499.900001n V_low
+ 500.000000n V_low
+ 500.000001n V_hig
+ 500.100000n V_hig
+ 500.100001n V_hig
+ 500.200000n V_hig
+ 500.200001n V_hig
+ 500.300000n V_hig
+ 500.300001n V_hig
+ 500.400000n V_hig
+ 500.400001n V_hig
+ 500.500000n V_hig
+ 500.500001n V_hig
+ 500.600000n V_hig
+ 500.600001n V_hig
+ 500.700000n V_hig
+ 500.700001n V_hig
+ 500.800000n V_hig
+ 500.800001n V_hig
+ 500.900000n V_hig
+ 500.900001n V_hig
+ 501.000000n V_hig
+ 501.000001n V_low
+ 501.100000n V_low
+ 501.100001n V_low
+ 501.200000n V_low
+ 501.200001n V_low
+ 501.300000n V_low
+ 501.300001n V_low
+ 501.400000n V_low
+ 501.400001n V_low
+ 501.500000n V_low
+ 501.500001n V_low
+ 501.600000n V_low
+ 501.600001n V_low
+ 501.700000n V_low
+ 501.700001n V_low
+ 501.800000n V_low
+ 501.800001n V_low
+ 501.900000n V_low
+ 501.900001n V_low
+ 502.000000n V_low
+ 502.000001n V_low
+ 502.100000n V_low
+ 502.100001n V_low
+ 502.200000n V_low
+ 502.200001n V_low
+ 502.300000n V_low
+ 502.300001n V_low
+ 502.400000n V_low
+ 502.400001n V_low
+ 502.500000n V_low
+ 502.500001n V_low
+ 502.600000n V_low
+ 502.600001n V_low
+ 502.700000n V_low
+ 502.700001n V_low
+ 502.800000n V_low
+ 502.800001n V_low
+ 502.900000n V_low
+ 502.900001n V_low
+ 503.000000n V_low
+ 503.000001n V_hig
+ 503.100000n V_hig
+ 503.100001n V_hig
+ 503.200000n V_hig
+ 503.200001n V_hig
+ 503.300000n V_hig
+ 503.300001n V_hig
+ 503.400000n V_hig
+ 503.400001n V_hig
+ 503.500000n V_hig
+ 503.500001n V_hig
+ 503.600000n V_hig
+ 503.600001n V_hig
+ 503.700000n V_hig
+ 503.700001n V_hig
+ 503.800000n V_hig
+ 503.800001n V_hig
+ 503.900000n V_hig
+ 503.900001n V_hig
+ 504.000000n V_hig
+ 504.000001n V_low
+ 504.100000n V_low
+ 504.100001n V_low
+ 504.200000n V_low
+ 504.200001n V_low
+ 504.300000n V_low
+ 504.300001n V_low
+ 504.400000n V_low
+ 504.400001n V_low
+ 504.500000n V_low
+ 504.500001n V_low
+ 504.600000n V_low
+ 504.600001n V_low
+ 504.700000n V_low
+ 504.700001n V_low
+ 504.800000n V_low
+ 504.800001n V_low
+ 504.900000n V_low
+ 504.900001n V_low
+ 505.000000n V_low
+ 505.000001n V_hig
+ 505.100000n V_hig
+ 505.100001n V_hig
+ 505.200000n V_hig
+ 505.200001n V_hig
+ 505.300000n V_hig
+ 505.300001n V_hig
+ 505.400000n V_hig
+ 505.400001n V_hig
+ 505.500000n V_hig
+ 505.500001n V_hig
+ 505.600000n V_hig
+ 505.600001n V_hig
+ 505.700000n V_hig
+ 505.700001n V_hig
+ 505.800000n V_hig
+ 505.800001n V_hig
+ 505.900000n V_hig
+ 505.900001n V_hig
+ 506.000000n V_hig
+ 506.000001n V_hig
+ 506.100000n V_hig
+ 506.100001n V_hig
+ 506.200000n V_hig
+ 506.200001n V_hig
+ 506.300000n V_hig
+ 506.300001n V_hig
+ 506.400000n V_hig
+ 506.400001n V_hig
+ 506.500000n V_hig
+ 506.500001n V_hig
+ 506.600000n V_hig
+ 506.600001n V_hig
+ 506.700000n V_hig
+ 506.700001n V_hig
+ 506.800000n V_hig
+ 506.800001n V_hig
+ 506.900000n V_hig
+ 506.900001n V_hig
+ 507.000000n V_hig
+ 507.000001n V_hig
+ 507.100000n V_hig
+ 507.100001n V_hig
+ 507.200000n V_hig
+ 507.200001n V_hig
+ 507.300000n V_hig
+ 507.300001n V_hig
+ 507.400000n V_hig
+ 507.400001n V_hig
+ 507.500000n V_hig
+ 507.500001n V_hig
+ 507.600000n V_hig
+ 507.600001n V_hig
+ 507.700000n V_hig
+ 507.700001n V_hig
+ 507.800000n V_hig
+ 507.800001n V_hig
+ 507.900000n V_hig
+ 507.900001n V_hig
+ 508.000000n V_hig
+ 508.000001n V_low
+ 508.100000n V_low
+ 508.100001n V_low
+ 508.200000n V_low
+ 508.200001n V_low
+ 508.300000n V_low
+ 508.300001n V_low
+ 508.400000n V_low
+ 508.400001n V_low
+ 508.500000n V_low
+ 508.500001n V_low
+ 508.600000n V_low
+ 508.600001n V_low
+ 508.700000n V_low
+ 508.700001n V_low
+ 508.800000n V_low
+ 508.800001n V_low
+ 508.900000n V_low
+ 508.900001n V_low
+ 509.000000n V_low
+ 509.000001n V_hig
+ 509.100000n V_hig
+ 509.100001n V_hig
+ 509.200000n V_hig
+ 509.200001n V_hig
+ 509.300000n V_hig
+ 509.300001n V_hig
+ 509.400000n V_hig
+ 509.400001n V_hig
+ 509.500000n V_hig
+ 509.500001n V_hig
+ 509.600000n V_hig
+ 509.600001n V_hig
+ 509.700000n V_hig
+ 509.700001n V_hig
+ 509.800000n V_hig
+ 509.800001n V_hig
+ 509.900000n V_hig
+ 509.900001n V_hig
+ 510.000000n V_hig
+ 510.000001n V_low
+ 510.100000n V_low
+ 510.100001n V_low
+ 510.200000n V_low
+ 510.200001n V_low
+ 510.300000n V_low
+ 510.300001n V_low
+ 510.400000n V_low
+ 510.400001n V_low
+ 510.500000n V_low
+ 510.500001n V_low
+ 510.600000n V_low
+ 510.600001n V_low
+ 510.700000n V_low
+ 510.700001n V_low
+ 510.800000n V_low
+ 510.800001n V_low
+ 510.900000n V_low
+ 510.900001n V_low
+ 511.000000n V_low
+ 511.000001n V_low
+ 511.100000n V_low
+ 511.100001n V_low
+ 511.200000n V_low
+ 511.200001n V_low
+ 511.300000n V_low
+ 511.300001n V_low
+ 511.400000n V_low
+ 511.400001n V_low
+ 511.500000n V_low
+ 511.500001n V_low
+ 511.600000n V_low
+ 511.600001n V_low
+ 511.700000n V_low
+ 511.700001n V_low
+ 511.800000n V_low
+ 511.800001n V_low
+ 511.900000n V_low
+ 511.900001n V_low
+ 512.000000n V_low
+ 512.000001n V_hig
+ 512.100000n V_hig
+ 512.100001n V_hig
+ 512.200000n V_hig
+ 512.200001n V_hig
+ 512.300000n V_hig
+ 512.300001n V_hig
+ 512.400000n V_hig
+ 512.400001n V_hig
+ 512.500000n V_hig
+ 512.500001n V_hig
+ 512.600000n V_hig
+ 512.600001n V_hig
+ 512.700000n V_hig
+ 512.700001n V_hig
+ 512.800000n V_hig
+ 512.800001n V_hig
+ 512.900000n V_hig
+ 512.900001n V_hig
+ 513.000000n V_hig
+ 513.000001n V_low
+ 513.100000n V_low
+ 513.100001n V_low
+ 513.200000n V_low
+ 513.200001n V_low
+ 513.300000n V_low
+ 513.300001n V_low
+ 513.400000n V_low
+ 513.400001n V_low
+ 513.500000n V_low
+ 513.500001n V_low
+ 513.600000n V_low
+ 513.600001n V_low
+ 513.700000n V_low
+ 513.700001n V_low
+ 513.800000n V_low
+ 513.800001n V_low
+ 513.900000n V_low
+ 513.900001n V_low
+ 514.000000n V_low
+ 514.000001n V_low
+ 514.100000n V_low
+ 514.100001n V_low
+ 514.200000n V_low
+ 514.200001n V_low
+ 514.300000n V_low
+ 514.300001n V_low
+ 514.400000n V_low
+ 514.400001n V_low
+ 514.500000n V_low
+ 514.500001n V_low
+ 514.600000n V_low
+ 514.600001n V_low
+ 514.700000n V_low
+ 514.700001n V_low
+ 514.800000n V_low
+ 514.800001n V_low
+ 514.900000n V_low
+ 514.900001n V_low
+ 515.000000n V_low
+ 515.000001n V_hig
+ 515.100000n V_hig
+ 515.100001n V_hig
+ 515.200000n V_hig
+ 515.200001n V_hig
+ 515.300000n V_hig
+ 515.300001n V_hig
+ 515.400000n V_hig
+ 515.400001n V_hig
+ 515.500000n V_hig
+ 515.500001n V_hig
+ 515.600000n V_hig
+ 515.600001n V_hig
+ 515.700000n V_hig
+ 515.700001n V_hig
+ 515.800000n V_hig
+ 515.800001n V_hig
+ 515.900000n V_hig
+ 515.900001n V_hig
+ 516.000000n V_hig
+ 516.000001n V_hig
+ 516.100000n V_hig
+ 516.100001n V_hig
+ 516.200000n V_hig
+ 516.200001n V_hig
+ 516.300000n V_hig
+ 516.300001n V_hig
+ 516.400000n V_hig
+ 516.400001n V_hig
+ 516.500000n V_hig
+ 516.500001n V_hig
+ 516.600000n V_hig
+ 516.600001n V_hig
+ 516.700000n V_hig
+ 516.700001n V_hig
+ 516.800000n V_hig
+ 516.800001n V_hig
+ 516.900000n V_hig
+ 516.900001n V_hig
+ 517.000000n V_hig
+ 517.000001n V_hig
+ 517.100000n V_hig
+ 517.100001n V_hig
+ 517.200000n V_hig
+ 517.200001n V_hig
+ 517.300000n V_hig
+ 517.300001n V_hig
+ 517.400000n V_hig
+ 517.400001n V_hig
+ 517.500000n V_hig
+ 517.500001n V_hig
+ 517.600000n V_hig
+ 517.600001n V_hig
+ 517.700000n V_hig
+ 517.700001n V_hig
+ 517.800000n V_hig
+ 517.800001n V_hig
+ 517.900000n V_hig
+ 517.900001n V_hig
+ 518.000000n V_hig
+ 518.000001n V_low
+ 518.100000n V_low
+ 518.100001n V_low
+ 518.200000n V_low
+ 518.200001n V_low
+ 518.300000n V_low
+ 518.300001n V_low
+ 518.400000n V_low
+ 518.400001n V_low
+ 518.500000n V_low
+ 518.500001n V_low
+ 518.600000n V_low
+ 518.600001n V_low
+ 518.700000n V_low
+ 518.700001n V_low
+ 518.800000n V_low
+ 518.800001n V_low
+ 518.900000n V_low
+ 518.900001n V_low
+ 519.000000n V_low
+ 519.000001n V_hig
+ 519.100000n V_hig
+ 519.100001n V_hig
+ 519.200000n V_hig
+ 519.200001n V_hig
+ 519.300000n V_hig
+ 519.300001n V_hig
+ 519.400000n V_hig
+ 519.400001n V_hig
+ 519.500000n V_hig
+ 519.500001n V_hig
+ 519.600000n V_hig
+ 519.600001n V_hig
+ 519.700000n V_hig
+ 519.700001n V_hig
+ 519.800000n V_hig
+ 519.800001n V_hig
+ 519.900000n V_hig
+ 519.900001n V_hig
+ 520.000000n V_hig
+ 520.000001n V_hig
+ 520.100000n V_hig
+ 520.100001n V_hig
+ 520.200000n V_hig
+ 520.200001n V_hig
+ 520.300000n V_hig
+ 520.300001n V_hig
+ 520.400000n V_hig
+ 520.400001n V_hig
+ 520.500000n V_hig
+ 520.500001n V_hig
+ 520.600000n V_hig
+ 520.600001n V_hig
+ 520.700000n V_hig
+ 520.700001n V_hig
+ 520.800000n V_hig
+ 520.800001n V_hig
+ 520.900000n V_hig
+ 520.900001n V_hig
+ 521.000000n V_hig
+ 521.000001n V_hig
+ 521.100000n V_hig
+ 521.100001n V_hig
+ 521.200000n V_hig
+ 521.200001n V_hig
+ 521.300000n V_hig
+ 521.300001n V_hig
+ 521.400000n V_hig
+ 521.400001n V_hig
+ 521.500000n V_hig
+ 521.500001n V_hig
+ 521.600000n V_hig
+ 521.600001n V_hig
+ 521.700000n V_hig
+ 521.700001n V_hig
+ 521.800000n V_hig
+ 521.800001n V_hig
+ 521.900000n V_hig
+ 521.900001n V_hig
+ 522.000000n V_hig
+ 522.000001n V_hig
+ 522.100000n V_hig
+ 522.100001n V_hig
+ 522.200000n V_hig
+ 522.200001n V_hig
+ 522.300000n V_hig
+ 522.300001n V_hig
+ 522.400000n V_hig
+ 522.400001n V_hig
+ 522.500000n V_hig
+ 522.500001n V_hig
+ 522.600000n V_hig
+ 522.600001n V_hig
+ 522.700000n V_hig
+ 522.700001n V_hig
+ 522.800000n V_hig
+ 522.800001n V_hig
+ 522.900000n V_hig
+ 522.900001n V_hig
+ 523.000000n V_hig
+ 523.000001n V_hig
+ 523.100000n V_hig
+ 523.100001n V_hig
+ 523.200000n V_hig
+ 523.200001n V_hig
+ 523.300000n V_hig
+ 523.300001n V_hig
+ 523.400000n V_hig
+ 523.400001n V_hig
+ 523.500000n V_hig
+ 523.500001n V_hig
+ 523.600000n V_hig
+ 523.600001n V_hig
+ 523.700000n V_hig
+ 523.700001n V_hig
+ 523.800000n V_hig
+ 523.800001n V_hig
+ 523.900000n V_hig
+ 523.900001n V_hig
+ 524.000000n V_hig
+ 524.000001n V_low
+ 524.100000n V_low
+ 524.100001n V_low
+ 524.200000n V_low
+ 524.200001n V_low
+ 524.300000n V_low
+ 524.300001n V_low
+ 524.400000n V_low
+ 524.400001n V_low
+ 524.500000n V_low
+ 524.500001n V_low
+ 524.600000n V_low
+ 524.600001n V_low
+ 524.700000n V_low
+ 524.700001n V_low
+ 524.800000n V_low
+ 524.800001n V_low
+ 524.900000n V_low
+ 524.900001n V_low
+ 525.000000n V_low
+ 525.000001n V_low
+ 525.100000n V_low
+ 525.100001n V_low
+ 525.200000n V_low
+ 525.200001n V_low
+ 525.300000n V_low
+ 525.300001n V_low
+ 525.400000n V_low
+ 525.400001n V_low
+ 525.500000n V_low
+ 525.500001n V_low
+ 525.600000n V_low
+ 525.600001n V_low
+ 525.700000n V_low
+ 525.700001n V_low
+ 525.800000n V_low
+ 525.800001n V_low
+ 525.900000n V_low
+ 525.900001n V_low
+ 526.000000n V_low
+ 526.000001n V_hig
+ 526.100000n V_hig
+ 526.100001n V_hig
+ 526.200000n V_hig
+ 526.200001n V_hig
+ 526.300000n V_hig
+ 526.300001n V_hig
+ 526.400000n V_hig
+ 526.400001n V_hig
+ 526.500000n V_hig
+ 526.500001n V_hig
+ 526.600000n V_hig
+ 526.600001n V_hig
+ 526.700000n V_hig
+ 526.700001n V_hig
+ 526.800000n V_hig
+ 526.800001n V_hig
+ 526.900000n V_hig
+ 526.900001n V_hig
+ 527.000000n V_hig
+ 527.000001n V_hig
+ 527.100000n V_hig
+ 527.100001n V_hig
+ 527.200000n V_hig
+ 527.200001n V_hig
+ 527.300000n V_hig
+ 527.300001n V_hig
+ 527.400000n V_hig
+ 527.400001n V_hig
+ 527.500000n V_hig
+ 527.500001n V_hig
+ 527.600000n V_hig
+ 527.600001n V_hig
+ 527.700000n V_hig
+ 527.700001n V_hig
+ 527.800000n V_hig
+ 527.800001n V_hig
+ 527.900000n V_hig
+ 527.900001n V_hig
+ 528.000000n V_hig
+ 528.000001n V_low
+ 528.100000n V_low
+ 528.100001n V_low
+ 528.200000n V_low
+ 528.200001n V_low
+ 528.300000n V_low
+ 528.300001n V_low
+ 528.400000n V_low
+ 528.400001n V_low
+ 528.500000n V_low
+ 528.500001n V_low
+ 528.600000n V_low
+ 528.600001n V_low
+ 528.700000n V_low
+ 528.700001n V_low
+ 528.800000n V_low
+ 528.800001n V_low
+ 528.900000n V_low
+ 528.900001n V_low
+ 529.000000n V_low
+ 529.000001n V_low
+ 529.100000n V_low
+ 529.100001n V_low
+ 529.200000n V_low
+ 529.200001n V_low
+ 529.300000n V_low
+ 529.300001n V_low
+ 529.400000n V_low
+ 529.400001n V_low
+ 529.500000n V_low
+ 529.500001n V_low
+ 529.600000n V_low
+ 529.600001n V_low
+ 529.700000n V_low
+ 529.700001n V_low
+ 529.800000n V_low
+ 529.800001n V_low
+ 529.900000n V_low
+ 529.900001n V_low
+ 530.000000n V_low
+ 530.000001n V_low
+ 530.100000n V_low
+ 530.100001n V_low
+ 530.200000n V_low
+ 530.200001n V_low
+ 530.300000n V_low
+ 530.300001n V_low
+ 530.400000n V_low
+ 530.400001n V_low
+ 530.500000n V_low
+ 530.500001n V_low
+ 530.600000n V_low
+ 530.600001n V_low
+ 530.700000n V_low
+ 530.700001n V_low
+ 530.800000n V_low
+ 530.800001n V_low
+ 530.900000n V_low
+ 530.900001n V_low
+ 531.000000n V_low
+ 531.000001n V_low
+ 531.100000n V_low
+ 531.100001n V_low
+ 531.200000n V_low
+ 531.200001n V_low
+ 531.300000n V_low
+ 531.300001n V_low
+ 531.400000n V_low
+ 531.400001n V_low
+ 531.500000n V_low
+ 531.500001n V_low
+ 531.600000n V_low
+ 531.600001n V_low
+ 531.700000n V_low
+ 531.700001n V_low
+ 531.800000n V_low
+ 531.800001n V_low
+ 531.900000n V_low
+ 531.900001n V_low
+ 532.000000n V_low
+ 532.000001n V_hig
+ 532.100000n V_hig
+ 532.100001n V_hig
+ 532.200000n V_hig
+ 532.200001n V_hig
+ 532.300000n V_hig
+ 532.300001n V_hig
+ 532.400000n V_hig
+ 532.400001n V_hig
+ 532.500000n V_hig
+ 532.500001n V_hig
+ 532.600000n V_hig
+ 532.600001n V_hig
+ 532.700000n V_hig
+ 532.700001n V_hig
+ 532.800000n V_hig
+ 532.800001n V_hig
+ 532.900000n V_hig
+ 532.900001n V_hig
+ 533.000000n V_hig
+ 533.000001n V_hig
+ 533.100000n V_hig
+ 533.100001n V_hig
+ 533.200000n V_hig
+ 533.200001n V_hig
+ 533.300000n V_hig
+ 533.300001n V_hig
+ 533.400000n V_hig
+ 533.400001n V_hig
+ 533.500000n V_hig
+ 533.500001n V_hig
+ 533.600000n V_hig
+ 533.600001n V_hig
+ 533.700000n V_hig
+ 533.700001n V_hig
+ 533.800000n V_hig
+ 533.800001n V_hig
+ 533.900000n V_hig
+ 533.900001n V_hig
+ 534.000000n V_hig
+ 534.000001n V_hig
+ 534.100000n V_hig
+ 534.100001n V_hig
+ 534.200000n V_hig
+ 534.200001n V_hig
+ 534.300000n V_hig
+ 534.300001n V_hig
+ 534.400000n V_hig
+ 534.400001n V_hig
+ 534.500000n V_hig
+ 534.500001n V_hig
+ 534.600000n V_hig
+ 534.600001n V_hig
+ 534.700000n V_hig
+ 534.700001n V_hig
+ 534.800000n V_hig
+ 534.800001n V_hig
+ 534.900000n V_hig
+ 534.900001n V_hig
+ 535.000000n V_hig
+ 535.000001n V_low
+ 535.100000n V_low
+ 535.100001n V_low
+ 535.200000n V_low
+ 535.200001n V_low
+ 535.300000n V_low
+ 535.300001n V_low
+ 535.400000n V_low
+ 535.400001n V_low
+ 535.500000n V_low
+ 535.500001n V_low
+ 535.600000n V_low
+ 535.600001n V_low
+ 535.700000n V_low
+ 535.700001n V_low
+ 535.800000n V_low
+ 535.800001n V_low
+ 535.900000n V_low
+ 535.900001n V_low
+ 536.000000n V_low
+ 536.000001n V_hig
+ 536.100000n V_hig
+ 536.100001n V_hig
+ 536.200000n V_hig
+ 536.200001n V_hig
+ 536.300000n V_hig
+ 536.300001n V_hig
+ 536.400000n V_hig
+ 536.400001n V_hig
+ 536.500000n V_hig
+ 536.500001n V_hig
+ 536.600000n V_hig
+ 536.600001n V_hig
+ 536.700000n V_hig
+ 536.700001n V_hig
+ 536.800000n V_hig
+ 536.800001n V_hig
+ 536.900000n V_hig
+ 536.900001n V_hig
+ 537.000000n V_hig
+ 537.000001n V_low
+ 537.100000n V_low
+ 537.100001n V_low
+ 537.200000n V_low
+ 537.200001n V_low
+ 537.300000n V_low
+ 537.300001n V_low
+ 537.400000n V_low
+ 537.400001n V_low
+ 537.500000n V_low
+ 537.500001n V_low
+ 537.600000n V_low
+ 537.600001n V_low
+ 537.700000n V_low
+ 537.700001n V_low
+ 537.800000n V_low
+ 537.800001n V_low
+ 537.900000n V_low
+ 537.900001n V_low
+ 538.000000n V_low
+ 538.000001n V_low
+ 538.100000n V_low
+ 538.100001n V_low
+ 538.200000n V_low
+ 538.200001n V_low
+ 538.300000n V_low
+ 538.300001n V_low
+ 538.400000n V_low
+ 538.400001n V_low
+ 538.500000n V_low
+ 538.500001n V_low
+ 538.600000n V_low
+ 538.600001n V_low
+ 538.700000n V_low
+ 538.700001n V_low
+ 538.800000n V_low
+ 538.800001n V_low
+ 538.900000n V_low
+ 538.900001n V_low
+ 539.000000n V_low
+ 539.000001n V_low
+ 539.100000n V_low
+ 539.100001n V_low
+ 539.200000n V_low
+ 539.200001n V_low
+ 539.300000n V_low
+ 539.300001n V_low
+ 539.400000n V_low
+ 539.400001n V_low
+ 539.500000n V_low
+ 539.500001n V_low
+ 539.600000n V_low
+ 539.600001n V_low
+ 539.700000n V_low
+ 539.700001n V_low
+ 539.800000n V_low
+ 539.800001n V_low
+ 539.900000n V_low
+ 539.900001n V_low
+ 540.000000n V_low
+ 540.000001n V_hig
+ 540.100000n V_hig
+ 540.100001n V_hig
+ 540.200000n V_hig
+ 540.200001n V_hig
+ 540.300000n V_hig
+ 540.300001n V_hig
+ 540.400000n V_hig
+ 540.400001n V_hig
+ 540.500000n V_hig
+ 540.500001n V_hig
+ 540.600000n V_hig
+ 540.600001n V_hig
+ 540.700000n V_hig
+ 540.700001n V_hig
+ 540.800000n V_hig
+ 540.800001n V_hig
+ 540.900000n V_hig
+ 540.900001n V_hig
+ 541.000000n V_hig
+ 541.000001n V_low
+ 541.100000n V_low
+ 541.100001n V_low
+ 541.200000n V_low
+ 541.200001n V_low
+ 541.300000n V_low
+ 541.300001n V_low
+ 541.400000n V_low
+ 541.400001n V_low
+ 541.500000n V_low
+ 541.500001n V_low
+ 541.600000n V_low
+ 541.600001n V_low
+ 541.700000n V_low
+ 541.700001n V_low
+ 541.800000n V_low
+ 541.800001n V_low
+ 541.900000n V_low
+ 541.900001n V_low
+ 542.000000n V_low
+ 542.000001n V_hig
+ 542.100000n V_hig
+ 542.100001n V_hig
+ 542.200000n V_hig
+ 542.200001n V_hig
+ 542.300000n V_hig
+ 542.300001n V_hig
+ 542.400000n V_hig
+ 542.400001n V_hig
+ 542.500000n V_hig
+ 542.500001n V_hig
+ 542.600000n V_hig
+ 542.600001n V_hig
+ 542.700000n V_hig
+ 542.700001n V_hig
+ 542.800000n V_hig
+ 542.800001n V_hig
+ 542.900000n V_hig
+ 542.900001n V_hig
+ 543.000000n V_hig
+ 543.000001n V_low
+ 543.100000n V_low
+ 543.100001n V_low
+ 543.200000n V_low
+ 543.200001n V_low
+ 543.300000n V_low
+ 543.300001n V_low
+ 543.400000n V_low
+ 543.400001n V_low
+ 543.500000n V_low
+ 543.500001n V_low
+ 543.600000n V_low
+ 543.600001n V_low
+ 543.700000n V_low
+ 543.700001n V_low
+ 543.800000n V_low
+ 543.800001n V_low
+ 543.900000n V_low
+ 543.900001n V_low
+ 544.000000n V_low
+ 544.000001n V_hig
+ 544.100000n V_hig
+ 544.100001n V_hig
+ 544.200000n V_hig
+ 544.200001n V_hig
+ 544.300000n V_hig
+ 544.300001n V_hig
+ 544.400000n V_hig
+ 544.400001n V_hig
+ 544.500000n V_hig
+ 544.500001n V_hig
+ 544.600000n V_hig
+ 544.600001n V_hig
+ 544.700000n V_hig
+ 544.700001n V_hig
+ 544.800000n V_hig
+ 544.800001n V_hig
+ 544.900000n V_hig
+ 544.900001n V_hig
+ 545.000000n V_hig
+ 545.000001n V_hig
+ 545.100000n V_hig
+ 545.100001n V_hig
+ 545.200000n V_hig
+ 545.200001n V_hig
+ 545.300000n V_hig
+ 545.300001n V_hig
+ 545.400000n V_hig
+ 545.400001n V_hig
+ 545.500000n V_hig
+ 545.500001n V_hig
+ 545.600000n V_hig
+ 545.600001n V_hig
+ 545.700000n V_hig
+ 545.700001n V_hig
+ 545.800000n V_hig
+ 545.800001n V_hig
+ 545.900000n V_hig
+ 545.900001n V_hig
+ 546.000000n V_hig
+ 546.000001n V_low
+ 546.100000n V_low
+ 546.100001n V_low
+ 546.200000n V_low
+ 546.200001n V_low
+ 546.300000n V_low
+ 546.300001n V_low
+ 546.400000n V_low
+ 546.400001n V_low
+ 546.500000n V_low
+ 546.500001n V_low
+ 546.600000n V_low
+ 546.600001n V_low
+ 546.700000n V_low
+ 546.700001n V_low
+ 546.800000n V_low
+ 546.800001n V_low
+ 546.900000n V_low
+ 546.900001n V_low
+ 547.000000n V_low
+ 547.000001n V_low
+ 547.100000n V_low
+ 547.100001n V_low
+ 547.200000n V_low
+ 547.200001n V_low
+ 547.300000n V_low
+ 547.300001n V_low
+ 547.400000n V_low
+ 547.400001n V_low
+ 547.500000n V_low
+ 547.500001n V_low
+ 547.600000n V_low
+ 547.600001n V_low
+ 547.700000n V_low
+ 547.700001n V_low
+ 547.800000n V_low
+ 547.800001n V_low
+ 547.900000n V_low
+ 547.900001n V_low
+ 548.000000n V_low
+ 548.000001n V_low
+ 548.100000n V_low
+ 548.100001n V_low
+ 548.200000n V_low
+ 548.200001n V_low
+ 548.300000n V_low
+ 548.300001n V_low
+ 548.400000n V_low
+ 548.400001n V_low
+ 548.500000n V_low
+ 548.500001n V_low
+ 548.600000n V_low
+ 548.600001n V_low
+ 548.700000n V_low
+ 548.700001n V_low
+ 548.800000n V_low
+ 548.800001n V_low
+ 548.900000n V_low
+ 548.900001n V_low
+ 549.000000n V_low
+ 549.000001n V_low
+ 549.100000n V_low
+ 549.100001n V_low
+ 549.200000n V_low
+ 549.200001n V_low
+ 549.300000n V_low
+ 549.300001n V_low
+ 549.400000n V_low
+ 549.400001n V_low
+ 549.500000n V_low
+ 549.500001n V_low
+ 549.600000n V_low
+ 549.600001n V_low
+ 549.700000n V_low
+ 549.700001n V_low
+ 549.800000n V_low
+ 549.800001n V_low
+ 549.900000n V_low
+ 549.900001n V_low
+ 550.000000n V_low
+ 550.000001n V_low
+ 550.100000n V_low
+ 550.100001n V_low
+ 550.200000n V_low
+ 550.200001n V_low
+ 550.300000n V_low
+ 550.300001n V_low
+ 550.400000n V_low
+ 550.400001n V_low
+ 550.500000n V_low
+ 550.500001n V_low
+ 550.600000n V_low
+ 550.600001n V_low
+ 550.700000n V_low
+ 550.700001n V_low
+ 550.800000n V_low
+ 550.800001n V_low
+ 550.900000n V_low
+ 550.900001n V_low
+ 551.000000n V_low
+ 551.000001n V_low
+ 551.100000n V_low
+ 551.100001n V_low
+ 551.200000n V_low
+ 551.200001n V_low
+ 551.300000n V_low
+ 551.300001n V_low
+ 551.400000n V_low
+ 551.400001n V_low
+ 551.500000n V_low
+ 551.500001n V_low
+ 551.600000n V_low
+ 551.600001n V_low
+ 551.700000n V_low
+ 551.700001n V_low
+ 551.800000n V_low
+ 551.800001n V_low
+ 551.900000n V_low
+ 551.900001n V_low
+ 552.000000n V_low
+ 552.000001n V_low
+ 552.100000n V_low
+ 552.100001n V_low
+ 552.200000n V_low
+ 552.200001n V_low
+ 552.300000n V_low
+ 552.300001n V_low
+ 552.400000n V_low
+ 552.400001n V_low
+ 552.500000n V_low
+ 552.500001n V_low
+ 552.600000n V_low
+ 552.600001n V_low
+ 552.700000n V_low
+ 552.700001n V_low
+ 552.800000n V_low
+ 552.800001n V_low
+ 552.900000n V_low
+ 552.900001n V_low
+ 553.000000n V_low
+ 553.000001n V_hig
+ 553.100000n V_hig
+ 553.100001n V_hig
+ 553.200000n V_hig
+ 553.200001n V_hig
+ 553.300000n V_hig
+ 553.300001n V_hig
+ 553.400000n V_hig
+ 553.400001n V_hig
+ 553.500000n V_hig
+ 553.500001n V_hig
+ 553.600000n V_hig
+ 553.600001n V_hig
+ 553.700000n V_hig
+ 553.700001n V_hig
+ 553.800000n V_hig
+ 553.800001n V_hig
+ 553.900000n V_hig
+ 553.900001n V_hig
+ 554.000000n V_hig
+ 554.000001n V_low
+ 554.100000n V_low
+ 554.100001n V_low
+ 554.200000n V_low
+ 554.200001n V_low
+ 554.300000n V_low
+ 554.300001n V_low
+ 554.400000n V_low
+ 554.400001n V_low
+ 554.500000n V_low
+ 554.500001n V_low
+ 554.600000n V_low
+ 554.600001n V_low
+ 554.700000n V_low
+ 554.700001n V_low
+ 554.800000n V_low
+ 554.800001n V_low
+ 554.900000n V_low
+ 554.900001n V_low
+ 555.000000n V_low
+ 555.000001n V_hig
+ 555.100000n V_hig
+ 555.100001n V_hig
+ 555.200000n V_hig
+ 555.200001n V_hig
+ 555.300000n V_hig
+ 555.300001n V_hig
+ 555.400000n V_hig
+ 555.400001n V_hig
+ 555.500000n V_hig
+ 555.500001n V_hig
+ 555.600000n V_hig
+ 555.600001n V_hig
+ 555.700000n V_hig
+ 555.700001n V_hig
+ 555.800000n V_hig
+ 555.800001n V_hig
+ 555.900000n V_hig
+ 555.900001n V_hig
+ 556.000000n V_hig
+ 556.000001n V_low
+ 556.100000n V_low
+ 556.100001n V_low
+ 556.200000n V_low
+ 556.200001n V_low
+ 556.300000n V_low
+ 556.300001n V_low
+ 556.400000n V_low
+ 556.400001n V_low
+ 556.500000n V_low
+ 556.500001n V_low
+ 556.600000n V_low
+ 556.600001n V_low
+ 556.700000n V_low
+ 556.700001n V_low
+ 556.800000n V_low
+ 556.800001n V_low
+ 556.900000n V_low
+ 556.900001n V_low
+ 557.000000n V_low
+ 557.000001n V_hig
+ 557.100000n V_hig
+ 557.100001n V_hig
+ 557.200000n V_hig
+ 557.200001n V_hig
+ 557.300000n V_hig
+ 557.300001n V_hig
+ 557.400000n V_hig
+ 557.400001n V_hig
+ 557.500000n V_hig
+ 557.500001n V_hig
+ 557.600000n V_hig
+ 557.600001n V_hig
+ 557.700000n V_hig
+ 557.700001n V_hig
+ 557.800000n V_hig
+ 557.800001n V_hig
+ 557.900000n V_hig
+ 557.900001n V_hig
+ 558.000000n V_hig
+ 558.000001n V_hig
+ 558.100000n V_hig
+ 558.100001n V_hig
+ 558.200000n V_hig
+ 558.200001n V_hig
+ 558.300000n V_hig
+ 558.300001n V_hig
+ 558.400000n V_hig
+ 558.400001n V_hig
+ 558.500000n V_hig
+ 558.500001n V_hig
+ 558.600000n V_hig
+ 558.600001n V_hig
+ 558.700000n V_hig
+ 558.700001n V_hig
+ 558.800000n V_hig
+ 558.800001n V_hig
+ 558.900000n V_hig
+ 558.900001n V_hig
+ 559.000000n V_hig
+ 559.000001n V_low
+ 559.100000n V_low
+ 559.100001n V_low
+ 559.200000n V_low
+ 559.200001n V_low
+ 559.300000n V_low
+ 559.300001n V_low
+ 559.400000n V_low
+ 559.400001n V_low
+ 559.500000n V_low
+ 559.500001n V_low
+ 559.600000n V_low
+ 559.600001n V_low
+ 559.700000n V_low
+ 559.700001n V_low
+ 559.800000n V_low
+ 559.800001n V_low
+ 559.900000n V_low
+ 559.900001n V_low
+ 560.000000n V_low
+ 560.000001n V_hig
+ 560.100000n V_hig
+ 560.100001n V_hig
+ 560.200000n V_hig
+ 560.200001n V_hig
+ 560.300000n V_hig
+ 560.300001n V_hig
+ 560.400000n V_hig
+ 560.400001n V_hig
+ 560.500000n V_hig
+ 560.500001n V_hig
+ 560.600000n V_hig
+ 560.600001n V_hig
+ 560.700000n V_hig
+ 560.700001n V_hig
+ 560.800000n V_hig
+ 560.800001n V_hig
+ 560.900000n V_hig
+ 560.900001n V_hig
+ 561.000000n V_hig
+ 561.000001n V_hig
+ 561.100000n V_hig
+ 561.100001n V_hig
+ 561.200000n V_hig
+ 561.200001n V_hig
+ 561.300000n V_hig
+ 561.300001n V_hig
+ 561.400000n V_hig
+ 561.400001n V_hig
+ 561.500000n V_hig
+ 561.500001n V_hig
+ 561.600000n V_hig
+ 561.600001n V_hig
+ 561.700000n V_hig
+ 561.700001n V_hig
+ 561.800000n V_hig
+ 561.800001n V_hig
+ 561.900000n V_hig
+ 561.900001n V_hig
+ 562.000000n V_hig
+ 562.000001n V_low
+ 562.100000n V_low
+ 562.100001n V_low
+ 562.200000n V_low
+ 562.200001n V_low
+ 562.300000n V_low
+ 562.300001n V_low
+ 562.400000n V_low
+ 562.400001n V_low
+ 562.500000n V_low
+ 562.500001n V_low
+ 562.600000n V_low
+ 562.600001n V_low
+ 562.700000n V_low
+ 562.700001n V_low
+ 562.800000n V_low
+ 562.800001n V_low
+ 562.900000n V_low
+ 562.900001n V_low
+ 563.000000n V_low
+ 563.000001n V_low
+ 563.100000n V_low
+ 563.100001n V_low
+ 563.200000n V_low
+ 563.200001n V_low
+ 563.300000n V_low
+ 563.300001n V_low
+ 563.400000n V_low
+ 563.400001n V_low
+ 563.500000n V_low
+ 563.500001n V_low
+ 563.600000n V_low
+ 563.600001n V_low
+ 563.700000n V_low
+ 563.700001n V_low
+ 563.800000n V_low
+ 563.800001n V_low
+ 563.900000n V_low
+ 563.900001n V_low
+ 564.000000n V_low
+ 564.000001n V_low
+ 564.100000n V_low
+ 564.100001n V_low
+ 564.200000n V_low
+ 564.200001n V_low
+ 564.300000n V_low
+ 564.300001n V_low
+ 564.400000n V_low
+ 564.400001n V_low
+ 564.500000n V_low
+ 564.500001n V_low
+ 564.600000n V_low
+ 564.600001n V_low
+ 564.700000n V_low
+ 564.700001n V_low
+ 564.800000n V_low
+ 564.800001n V_low
+ 564.900000n V_low
+ 564.900001n V_low
+ 565.000000n V_low
+ 565.000001n V_hig
+ 565.100000n V_hig
+ 565.100001n V_hig
+ 565.200000n V_hig
+ 565.200001n V_hig
+ 565.300000n V_hig
+ 565.300001n V_hig
+ 565.400000n V_hig
+ 565.400001n V_hig
+ 565.500000n V_hig
+ 565.500001n V_hig
+ 565.600000n V_hig
+ 565.600001n V_hig
+ 565.700000n V_hig
+ 565.700001n V_hig
+ 565.800000n V_hig
+ 565.800001n V_hig
+ 565.900000n V_hig
+ 565.900001n V_hig
+ 566.000000n V_hig
+ 566.000001n V_low
+ 566.100000n V_low
+ 566.100001n V_low
+ 566.200000n V_low
+ 566.200001n V_low
+ 566.300000n V_low
+ 566.300001n V_low
+ 566.400000n V_low
+ 566.400001n V_low
+ 566.500000n V_low
+ 566.500001n V_low
+ 566.600000n V_low
+ 566.600001n V_low
+ 566.700000n V_low
+ 566.700001n V_low
+ 566.800000n V_low
+ 566.800001n V_low
+ 566.900000n V_low
+ 566.900001n V_low
+ 567.000000n V_low
+ 567.000001n V_low
+ 567.100000n V_low
+ 567.100001n V_low
+ 567.200000n V_low
+ 567.200001n V_low
+ 567.300000n V_low
+ 567.300001n V_low
+ 567.400000n V_low
+ 567.400001n V_low
+ 567.500000n V_low
+ 567.500001n V_low
+ 567.600000n V_low
+ 567.600001n V_low
+ 567.700000n V_low
+ 567.700001n V_low
+ 567.800000n V_low
+ 567.800001n V_low
+ 567.900000n V_low
+ 567.900001n V_low
+ 568.000000n V_low
+ 568.000001n V_low
+ 568.100000n V_low
+ 568.100001n V_low
+ 568.200000n V_low
+ 568.200001n V_low
+ 568.300000n V_low
+ 568.300001n V_low
+ 568.400000n V_low
+ 568.400001n V_low
+ 568.500000n V_low
+ 568.500001n V_low
+ 568.600000n V_low
+ 568.600001n V_low
+ 568.700000n V_low
+ 568.700001n V_low
+ 568.800000n V_low
+ 568.800001n V_low
+ 568.900000n V_low
+ 568.900001n V_low
+ 569.000000n V_low
+ 569.000001n V_low
+ 569.100000n V_low
+ 569.100001n V_low
+ 569.200000n V_low
+ 569.200001n V_low
+ 569.300000n V_low
+ 569.300001n V_low
+ 569.400000n V_low
+ 569.400001n V_low
+ 569.500000n V_low
+ 569.500001n V_low
+ 569.600000n V_low
+ 569.600001n V_low
+ 569.700000n V_low
+ 569.700001n V_low
+ 569.800000n V_low
+ 569.800001n V_low
+ 569.900000n V_low
+ 569.900001n V_low
+ 570.000000n V_low
+ 570.000001n V_hig
+ 570.100000n V_hig
+ 570.100001n V_hig
+ 570.200000n V_hig
+ 570.200001n V_hig
+ 570.300000n V_hig
+ 570.300001n V_hig
+ 570.400000n V_hig
+ 570.400001n V_hig
+ 570.500000n V_hig
+ 570.500001n V_hig
+ 570.600000n V_hig
+ 570.600001n V_hig
+ 570.700000n V_hig
+ 570.700001n V_hig
+ 570.800000n V_hig
+ 570.800001n V_hig
+ 570.900000n V_hig
+ 570.900001n V_hig
+ 571.000000n V_hig
+ 571.000001n V_hig
+ 571.100000n V_hig
+ 571.100001n V_hig
+ 571.200000n V_hig
+ 571.200001n V_hig
+ 571.300000n V_hig
+ 571.300001n V_hig
+ 571.400000n V_hig
+ 571.400001n V_hig
+ 571.500000n V_hig
+ 571.500001n V_hig
+ 571.600000n V_hig
+ 571.600001n V_hig
+ 571.700000n V_hig
+ 571.700001n V_hig
+ 571.800000n V_hig
+ 571.800001n V_hig
+ 571.900000n V_hig
+ 571.900001n V_hig
+ 572.000000n V_hig
+ 572.000001n V_hig
+ 572.100000n V_hig
+ 572.100001n V_hig
+ 572.200000n V_hig
+ 572.200001n V_hig
+ 572.300000n V_hig
+ 572.300001n V_hig
+ 572.400000n V_hig
+ 572.400001n V_hig
+ 572.500000n V_hig
+ 572.500001n V_hig
+ 572.600000n V_hig
+ 572.600001n V_hig
+ 572.700000n V_hig
+ 572.700001n V_hig
+ 572.800000n V_hig
+ 572.800001n V_hig
+ 572.900000n V_hig
+ 572.900001n V_hig
+ 573.000000n V_hig
+ 573.000001n V_low
+ 573.100000n V_low
+ 573.100001n V_low
+ 573.200000n V_low
+ 573.200001n V_low
+ 573.300000n V_low
+ 573.300001n V_low
+ 573.400000n V_low
+ 573.400001n V_low
+ 573.500000n V_low
+ 573.500001n V_low
+ 573.600000n V_low
+ 573.600001n V_low
+ 573.700000n V_low
+ 573.700001n V_low
+ 573.800000n V_low
+ 573.800001n V_low
+ 573.900000n V_low
+ 573.900001n V_low
+ 574.000000n V_low
+ 574.000001n V_low
+ 574.100000n V_low
+ 574.100001n V_low
+ 574.200000n V_low
+ 574.200001n V_low
+ 574.300000n V_low
+ 574.300001n V_low
+ 574.400000n V_low
+ 574.400001n V_low
+ 574.500000n V_low
+ 574.500001n V_low
+ 574.600000n V_low
+ 574.600001n V_low
+ 574.700000n V_low
+ 574.700001n V_low
+ 574.800000n V_low
+ 574.800001n V_low
+ 574.900000n V_low
+ 574.900001n V_low
+ 575.000000n V_low
+ 575.000001n V_hig
+ 575.100000n V_hig
+ 575.100001n V_hig
+ 575.200000n V_hig
+ 575.200001n V_hig
+ 575.300000n V_hig
+ 575.300001n V_hig
+ 575.400000n V_hig
+ 575.400001n V_hig
+ 575.500000n V_hig
+ 575.500001n V_hig
+ 575.600000n V_hig
+ 575.600001n V_hig
+ 575.700000n V_hig
+ 575.700001n V_hig
+ 575.800000n V_hig
+ 575.800001n V_hig
+ 575.900000n V_hig
+ 575.900001n V_hig
+ 576.000000n V_hig
+ 576.000001n V_hig
+ 576.100000n V_hig
+ 576.100001n V_hig
+ 576.200000n V_hig
+ 576.200001n V_hig
+ 576.300000n V_hig
+ 576.300001n V_hig
+ 576.400000n V_hig
+ 576.400001n V_hig
+ 576.500000n V_hig
+ 576.500001n V_hig
+ 576.600000n V_hig
+ 576.600001n V_hig
+ 576.700000n V_hig
+ 576.700001n V_hig
+ 576.800000n V_hig
+ 576.800001n V_hig
+ 576.900000n V_hig
+ 576.900001n V_hig
+ 577.000000n V_hig
+ 577.000001n V_low
+ 577.100000n V_low
+ 577.100001n V_low
+ 577.200000n V_low
+ 577.200001n V_low
+ 577.300000n V_low
+ 577.300001n V_low
+ 577.400000n V_low
+ 577.400001n V_low
+ 577.500000n V_low
+ 577.500001n V_low
+ 577.600000n V_low
+ 577.600001n V_low
+ 577.700000n V_low
+ 577.700001n V_low
+ 577.800000n V_low
+ 577.800001n V_low
+ 577.900000n V_low
+ 577.900001n V_low
+ 578.000000n V_low
+ 578.000001n V_low
+ 578.100000n V_low
+ 578.100001n V_low
+ 578.200000n V_low
+ 578.200001n V_low
+ 578.300000n V_low
+ 578.300001n V_low
+ 578.400000n V_low
+ 578.400001n V_low
+ 578.500000n V_low
+ 578.500001n V_low
+ 578.600000n V_low
+ 578.600001n V_low
+ 578.700000n V_low
+ 578.700001n V_low
+ 578.800000n V_low
+ 578.800001n V_low
+ 578.900000n V_low
+ 578.900001n V_low
+ 579.000000n V_low
+ 579.000001n V_hig
+ 579.100000n V_hig
+ 579.100001n V_hig
+ 579.200000n V_hig
+ 579.200001n V_hig
+ 579.300000n V_hig
+ 579.300001n V_hig
+ 579.400000n V_hig
+ 579.400001n V_hig
+ 579.500000n V_hig
+ 579.500001n V_hig
+ 579.600000n V_hig
+ 579.600001n V_hig
+ 579.700000n V_hig
+ 579.700001n V_hig
+ 579.800000n V_hig
+ 579.800001n V_hig
+ 579.900000n V_hig
+ 579.900001n V_hig
+ 580.000000n V_hig
+ 580.000001n V_low
+ 580.100000n V_low
+ 580.100001n V_low
+ 580.200000n V_low
+ 580.200001n V_low
+ 580.300000n V_low
+ 580.300001n V_low
+ 580.400000n V_low
+ 580.400001n V_low
+ 580.500000n V_low
+ 580.500001n V_low
+ 580.600000n V_low
+ 580.600001n V_low
+ 580.700000n V_low
+ 580.700001n V_low
+ 580.800000n V_low
+ 580.800001n V_low
+ 580.900000n V_low
+ 580.900001n V_low
+ 581.000000n V_low
+ 581.000001n V_hig
+ 581.100000n V_hig
+ 581.100001n V_hig
+ 581.200000n V_hig
+ 581.200001n V_hig
+ 581.300000n V_hig
+ 581.300001n V_hig
+ 581.400000n V_hig
+ 581.400001n V_hig
+ 581.500000n V_hig
+ 581.500001n V_hig
+ 581.600000n V_hig
+ 581.600001n V_hig
+ 581.700000n V_hig
+ 581.700001n V_hig
+ 581.800000n V_hig
+ 581.800001n V_hig
+ 581.900000n V_hig
+ 581.900001n V_hig
+ 582.000000n V_hig
+ 582.000001n V_hig
+ 582.100000n V_hig
+ 582.100001n V_hig
+ 582.200000n V_hig
+ 582.200001n V_hig
+ 582.300000n V_hig
+ 582.300001n V_hig
+ 582.400000n V_hig
+ 582.400001n V_hig
+ 582.500000n V_hig
+ 582.500001n V_hig
+ 582.600000n V_hig
+ 582.600001n V_hig
+ 582.700000n V_hig
+ 582.700001n V_hig
+ 582.800000n V_hig
+ 582.800001n V_hig
+ 582.900000n V_hig
+ 582.900001n V_hig
+ 583.000000n V_hig
+ 583.000001n V_hig
+ 583.100000n V_hig
+ 583.100001n V_hig
+ 583.200000n V_hig
+ 583.200001n V_hig
+ 583.300000n V_hig
+ 583.300001n V_hig
+ 583.400000n V_hig
+ 583.400001n V_hig
+ 583.500000n V_hig
+ 583.500001n V_hig
+ 583.600000n V_hig
+ 583.600001n V_hig
+ 583.700000n V_hig
+ 583.700001n V_hig
+ 583.800000n V_hig
+ 583.800001n V_hig
+ 583.900000n V_hig
+ 583.900001n V_hig
+ 584.000000n V_hig
+ 584.000001n V_hig
+ 584.100000n V_hig
+ 584.100001n V_hig
+ 584.200000n V_hig
+ 584.200001n V_hig
+ 584.300000n V_hig
+ 584.300001n V_hig
+ 584.400000n V_hig
+ 584.400001n V_hig
+ 584.500000n V_hig
+ 584.500001n V_hig
+ 584.600000n V_hig
+ 584.600001n V_hig
+ 584.700000n V_hig
+ 584.700001n V_hig
+ 584.800000n V_hig
+ 584.800001n V_hig
+ 584.900000n V_hig
+ 584.900001n V_hig
+ 585.000000n V_hig
+ 585.000001n V_hig
+ 585.100000n V_hig
+ 585.100001n V_hig
+ 585.200000n V_hig
+ 585.200001n V_hig
+ 585.300000n V_hig
+ 585.300001n V_hig
+ 585.400000n V_hig
+ 585.400001n V_hig
+ 585.500000n V_hig
+ 585.500001n V_hig
+ 585.600000n V_hig
+ 585.600001n V_hig
+ 585.700000n V_hig
+ 585.700001n V_hig
+ 585.800000n V_hig
+ 585.800001n V_hig
+ 585.900000n V_hig
+ 585.900001n V_hig
+ 586.000000n V_hig
+ 586.000001n V_hig
+ 586.100000n V_hig
+ 586.100001n V_hig
+ 586.200000n V_hig
+ 586.200001n V_hig
+ 586.300000n V_hig
+ 586.300001n V_hig
+ 586.400000n V_hig
+ 586.400001n V_hig
+ 586.500000n V_hig
+ 586.500001n V_hig
+ 586.600000n V_hig
+ 586.600001n V_hig
+ 586.700000n V_hig
+ 586.700001n V_hig
+ 586.800000n V_hig
+ 586.800001n V_hig
+ 586.900000n V_hig
+ 586.900001n V_hig
+ 587.000000n V_hig
+ 587.000001n V_low
+ 587.100000n V_low
+ 587.100001n V_low
+ 587.200000n V_low
+ 587.200001n V_low
+ 587.300000n V_low
+ 587.300001n V_low
+ 587.400000n V_low
+ 587.400001n V_low
+ 587.500000n V_low
+ 587.500001n V_low
+ 587.600000n V_low
+ 587.600001n V_low
+ 587.700000n V_low
+ 587.700001n V_low
+ 587.800000n V_low
+ 587.800001n V_low
+ 587.900000n V_low
+ 587.900001n V_low
+ 588.000000n V_low
+ 588.000001n V_hig
+ 588.100000n V_hig
+ 588.100001n V_hig
+ 588.200000n V_hig
+ 588.200001n V_hig
+ 588.300000n V_hig
+ 588.300001n V_hig
+ 588.400000n V_hig
+ 588.400001n V_hig
+ 588.500000n V_hig
+ 588.500001n V_hig
+ 588.600000n V_hig
+ 588.600001n V_hig
+ 588.700000n V_hig
+ 588.700001n V_hig
+ 588.800000n V_hig
+ 588.800001n V_hig
+ 588.900000n V_hig
+ 588.900001n V_hig
+ 589.000000n V_hig
+ 589.000001n V_hig
+ 589.100000n V_hig
+ 589.100001n V_hig
+ 589.200000n V_hig
+ 589.200001n V_hig
+ 589.300000n V_hig
+ 589.300001n V_hig
+ 589.400000n V_hig
+ 589.400001n V_hig
+ 589.500000n V_hig
+ 589.500001n V_hig
+ 589.600000n V_hig
+ 589.600001n V_hig
+ 589.700000n V_hig
+ 589.700001n V_hig
+ 589.800000n V_hig
+ 589.800001n V_hig
+ 589.900000n V_hig
+ 589.900001n V_hig
+ 590.000000n V_hig
+ 590.000001n V_low
+ 590.100000n V_low
+ 590.100001n V_low
+ 590.200000n V_low
+ 590.200001n V_low
+ 590.300000n V_low
+ 590.300001n V_low
+ 590.400000n V_low
+ 590.400001n V_low
+ 590.500000n V_low
+ 590.500001n V_low
+ 590.600000n V_low
+ 590.600001n V_low
+ 590.700000n V_low
+ 590.700001n V_low
+ 590.800000n V_low
+ 590.800001n V_low
+ 590.900000n V_low
+ 590.900001n V_low
+ 591.000000n V_low
+ 591.000001n V_hig
+ 591.100000n V_hig
+ 591.100001n V_hig
+ 591.200000n V_hig
+ 591.200001n V_hig
+ 591.300000n V_hig
+ 591.300001n V_hig
+ 591.400000n V_hig
+ 591.400001n V_hig
+ 591.500000n V_hig
+ 591.500001n V_hig
+ 591.600000n V_hig
+ 591.600001n V_hig
+ 591.700000n V_hig
+ 591.700001n V_hig
+ 591.800000n V_hig
+ 591.800001n V_hig
+ 591.900000n V_hig
+ 591.900001n V_hig
+ 592.000000n V_hig
+ 592.000001n V_low
+ 592.100000n V_low
+ 592.100001n V_low
+ 592.200000n V_low
+ 592.200001n V_low
+ 592.300000n V_low
+ 592.300001n V_low
+ 592.400000n V_low
+ 592.400001n V_low
+ 592.500000n V_low
+ 592.500001n V_low
+ 592.600000n V_low
+ 592.600001n V_low
+ 592.700000n V_low
+ 592.700001n V_low
+ 592.800000n V_low
+ 592.800001n V_low
+ 592.900000n V_low
+ 592.900001n V_low
+ 593.000000n V_low
+ 593.000001n V_low
+ 593.100000n V_low
+ 593.100001n V_low
+ 593.200000n V_low
+ 593.200001n V_low
+ 593.300000n V_low
+ 593.300001n V_low
+ 593.400000n V_low
+ 593.400001n V_low
+ 593.500000n V_low
+ 593.500001n V_low
+ 593.600000n V_low
+ 593.600001n V_low
+ 593.700000n V_low
+ 593.700001n V_low
+ 593.800000n V_low
+ 593.800001n V_low
+ 593.900000n V_low
+ 593.900001n V_low
+ 594.000000n V_low
+ 594.000001n V_hig
+ 594.100000n V_hig
+ 594.100001n V_hig
+ 594.200000n V_hig
+ 594.200001n V_hig
+ 594.300000n V_hig
+ 594.300001n V_hig
+ 594.400000n V_hig
+ 594.400001n V_hig
+ 594.500000n V_hig
+ 594.500001n V_hig
+ 594.600000n V_hig
+ 594.600001n V_hig
+ 594.700000n V_hig
+ 594.700001n V_hig
+ 594.800000n V_hig
+ 594.800001n V_hig
+ 594.900000n V_hig
+ 594.900001n V_hig
+ 595.000000n V_hig
+ 595.000001n V_hig
+ 595.100000n V_hig
+ 595.100001n V_hig
+ 595.200000n V_hig
+ 595.200001n V_hig
+ 595.300000n V_hig
+ 595.300001n V_hig
+ 595.400000n V_hig
+ 595.400001n V_hig
+ 595.500000n V_hig
+ 595.500001n V_hig
+ 595.600000n V_hig
+ 595.600001n V_hig
+ 595.700000n V_hig
+ 595.700001n V_hig
+ 595.800000n V_hig
+ 595.800001n V_hig
+ 595.900000n V_hig
+ 595.900001n V_hig
+ 596.000000n V_hig
+ 596.000001n V_hig
+ 596.100000n V_hig
+ 596.100001n V_hig
+ 596.200000n V_hig
+ 596.200001n V_hig
+ 596.300000n V_hig
+ 596.300001n V_hig
+ 596.400000n V_hig
+ 596.400001n V_hig
+ 596.500000n V_hig
+ 596.500001n V_hig
+ 596.600000n V_hig
+ 596.600001n V_hig
+ 596.700000n V_hig
+ 596.700001n V_hig
+ 596.800000n V_hig
+ 596.800001n V_hig
+ 596.900000n V_hig
+ 596.900001n V_hig
+ 597.000000n V_hig
+ 597.000001n V_low
+ 597.100000n V_low
+ 597.100001n V_low
+ 597.200000n V_low
+ 597.200001n V_low
+ 597.300000n V_low
+ 597.300001n V_low
+ 597.400000n V_low
+ 597.400001n V_low
+ 597.500000n V_low
+ 597.500001n V_low
+ 597.600000n V_low
+ 597.600001n V_low
+ 597.700000n V_low
+ 597.700001n V_low
+ 597.800000n V_low
+ 597.800001n V_low
+ 597.900000n V_low
+ 597.900001n V_low
+ 598.000000n V_low
+ 598.000001n V_hig
+ 598.100000n V_hig
+ 598.100001n V_hig
+ 598.200000n V_hig
+ 598.200001n V_hig
+ 598.300000n V_hig
+ 598.300001n V_hig
+ 598.400000n V_hig
+ 598.400001n V_hig
+ 598.500000n V_hig
+ 598.500001n V_hig
+ 598.600000n V_hig
+ 598.600001n V_hig
+ 598.700000n V_hig
+ 598.700001n V_hig
+ 598.800000n V_hig
+ 598.800001n V_hig
+ 598.900000n V_hig
+ 598.900001n V_hig
+ 599.000000n V_hig
+ 599.000001n V_low
+ 599.100000n V_low
+ 599.100001n V_low
+ 599.200000n V_low
+ 599.200001n V_low
+ 599.300000n V_low
+ 599.300001n V_low
+ 599.400000n V_low
+ 599.400001n V_low
+ 599.500000n V_low
+ 599.500001n V_low
+ 599.600000n V_low
+ 599.600001n V_low
+ 599.700000n V_low
+ 599.700001n V_low
+ 599.800000n V_low
+ 599.800001n V_low
+ 599.900000n V_low
+ 599.900001n V_low
+ 600.000000n V_low
+ 600.000001n V_hig
+ 600.100000n V_hig
+ 600.100001n V_hig
+ 600.200000n V_hig
+ 600.200001n V_hig
+ 600.300000n V_hig
+ 600.300001n V_hig
+ 600.400000n V_hig
+ 600.400001n V_hig
+ 600.500000n V_hig
+ 600.500001n V_hig
+ 600.600000n V_hig
+ 600.600001n V_hig
+ 600.700000n V_hig
+ 600.700001n V_hig
+ 600.800000n V_hig
+ 600.800001n V_hig
+ 600.900000n V_hig
+ 600.900001n V_hig
+ 601.000000n V_hig
+ 601.000001n V_hig
+ 601.100000n V_hig
+ 601.100001n V_hig
+ 601.200000n V_hig
+ 601.200001n V_hig
+ 601.300000n V_hig
+ 601.300001n V_hig
+ 601.400000n V_hig
+ 601.400001n V_hig
+ 601.500000n V_hig
+ 601.500001n V_hig
+ 601.600000n V_hig
+ 601.600001n V_hig
+ 601.700000n V_hig
+ 601.700001n V_hig
+ 601.800000n V_hig
+ 601.800001n V_hig
+ 601.900000n V_hig
+ 601.900001n V_hig
+ 602.000000n V_hig
+ 602.000001n V_hig
+ 602.100000n V_hig
+ 602.100001n V_hig
+ 602.200000n V_hig
+ 602.200001n V_hig
+ 602.300000n V_hig
+ 602.300001n V_hig
+ 602.400000n V_hig
+ 602.400001n V_hig
+ 602.500000n V_hig
+ 602.500001n V_hig
+ 602.600000n V_hig
+ 602.600001n V_hig
+ 602.700000n V_hig
+ 602.700001n V_hig
+ 602.800000n V_hig
+ 602.800001n V_hig
+ 602.900000n V_hig
+ 602.900001n V_hig
+ 603.000000n V_hig
+ 603.000001n V_low
+ 603.100000n V_low
+ 603.100001n V_low
+ 603.200000n V_low
+ 603.200001n V_low
+ 603.300000n V_low
+ 603.300001n V_low
+ 603.400000n V_low
+ 603.400001n V_low
+ 603.500000n V_low
+ 603.500001n V_low
+ 603.600000n V_low
+ 603.600001n V_low
+ 603.700000n V_low
+ 603.700001n V_low
+ 603.800000n V_low
+ 603.800001n V_low
+ 603.900000n V_low
+ 603.900001n V_low
+ 604.000000n V_low
+ 604.000001n V_low
+ 604.100000n V_low
+ 604.100001n V_low
+ 604.200000n V_low
+ 604.200001n V_low
+ 604.300000n V_low
+ 604.300001n V_low
+ 604.400000n V_low
+ 604.400001n V_low
+ 604.500000n V_low
+ 604.500001n V_low
+ 604.600000n V_low
+ 604.600001n V_low
+ 604.700000n V_low
+ 604.700001n V_low
+ 604.800000n V_low
+ 604.800001n V_low
+ 604.900000n V_low
+ 604.900001n V_low
+ 605.000000n V_low
+ 605.000001n V_hig
+ 605.100000n V_hig
+ 605.100001n V_hig
+ 605.200000n V_hig
+ 605.200001n V_hig
+ 605.300000n V_hig
+ 605.300001n V_hig
+ 605.400000n V_hig
+ 605.400001n V_hig
+ 605.500000n V_hig
+ 605.500001n V_hig
+ 605.600000n V_hig
+ 605.600001n V_hig
+ 605.700000n V_hig
+ 605.700001n V_hig
+ 605.800000n V_hig
+ 605.800001n V_hig
+ 605.900000n V_hig
+ 605.900001n V_hig
+ 606.000000n V_hig
+ 606.000001n V_low
+ 606.100000n V_low
+ 606.100001n V_low
+ 606.200000n V_low
+ 606.200001n V_low
+ 606.300000n V_low
+ 606.300001n V_low
+ 606.400000n V_low
+ 606.400001n V_low
+ 606.500000n V_low
+ 606.500001n V_low
+ 606.600000n V_low
+ 606.600001n V_low
+ 606.700000n V_low
+ 606.700001n V_low
+ 606.800000n V_low
+ 606.800001n V_low
+ 606.900000n V_low
+ 606.900001n V_low
+ 607.000000n V_low
+ 607.000001n V_hig
+ 607.100000n V_hig
+ 607.100001n V_hig
+ 607.200000n V_hig
+ 607.200001n V_hig
+ 607.300000n V_hig
+ 607.300001n V_hig
+ 607.400000n V_hig
+ 607.400001n V_hig
+ 607.500000n V_hig
+ 607.500001n V_hig
+ 607.600000n V_hig
+ 607.600001n V_hig
+ 607.700000n V_hig
+ 607.700001n V_hig
+ 607.800000n V_hig
+ 607.800001n V_hig
+ 607.900000n V_hig
+ 607.900001n V_hig
+ 608.000000n V_hig
+ 608.000001n V_hig
+ 608.100000n V_hig
+ 608.100001n V_hig
+ 608.200000n V_hig
+ 608.200001n V_hig
+ 608.300000n V_hig
+ 608.300001n V_hig
+ 608.400000n V_hig
+ 608.400001n V_hig
+ 608.500000n V_hig
+ 608.500001n V_hig
+ 608.600000n V_hig
+ 608.600001n V_hig
+ 608.700000n V_hig
+ 608.700001n V_hig
+ 608.800000n V_hig
+ 608.800001n V_hig
+ 608.900000n V_hig
+ 608.900001n V_hig
+ 609.000000n V_hig
+ 609.000001n V_low
+ 609.100000n V_low
+ 609.100001n V_low
+ 609.200000n V_low
+ 609.200001n V_low
+ 609.300000n V_low
+ 609.300001n V_low
+ 609.400000n V_low
+ 609.400001n V_low
+ 609.500000n V_low
+ 609.500001n V_low
+ 609.600000n V_low
+ 609.600001n V_low
+ 609.700000n V_low
+ 609.700001n V_low
+ 609.800000n V_low
+ 609.800001n V_low
+ 609.900000n V_low
+ 609.900001n V_low
+ 610.000000n V_low
+ 610.000001n V_hig
+ 610.100000n V_hig
+ 610.100001n V_hig
+ 610.200000n V_hig
+ 610.200001n V_hig
+ 610.300000n V_hig
+ 610.300001n V_hig
+ 610.400000n V_hig
+ 610.400001n V_hig
+ 610.500000n V_hig
+ 610.500001n V_hig
+ 610.600000n V_hig
+ 610.600001n V_hig
+ 610.700000n V_hig
+ 610.700001n V_hig
+ 610.800000n V_hig
+ 610.800001n V_hig
+ 610.900000n V_hig
+ 610.900001n V_hig
+ 611.000000n V_hig
+ 611.000001n V_hig
+ 611.100000n V_hig
+ 611.100001n V_hig
+ 611.200000n V_hig
+ 611.200001n V_hig
+ 611.300000n V_hig
+ 611.300001n V_hig
+ 611.400000n V_hig
+ 611.400001n V_hig
+ 611.500000n V_hig
+ 611.500001n V_hig
+ 611.600000n V_hig
+ 611.600001n V_hig
+ 611.700000n V_hig
+ 611.700001n V_hig
+ 611.800000n V_hig
+ 611.800001n V_hig
+ 611.900000n V_hig
+ 611.900001n V_hig
+ 612.000000n V_hig
+ 612.000001n V_low
+ 612.100000n V_low
+ 612.100001n V_low
+ 612.200000n V_low
+ 612.200001n V_low
+ 612.300000n V_low
+ 612.300001n V_low
+ 612.400000n V_low
+ 612.400001n V_low
+ 612.500000n V_low
+ 612.500001n V_low
+ 612.600000n V_low
+ 612.600001n V_low
+ 612.700000n V_low
+ 612.700001n V_low
+ 612.800000n V_low
+ 612.800001n V_low
+ 612.900000n V_low
+ 612.900001n V_low
+ 613.000000n V_low
+ 613.000001n V_low
+ 613.100000n V_low
+ 613.100001n V_low
+ 613.200000n V_low
+ 613.200001n V_low
+ 613.300000n V_low
+ 613.300001n V_low
+ 613.400000n V_low
+ 613.400001n V_low
+ 613.500000n V_low
+ 613.500001n V_low
+ 613.600000n V_low
+ 613.600001n V_low
+ 613.700000n V_low
+ 613.700001n V_low
+ 613.800000n V_low
+ 613.800001n V_low
+ 613.900000n V_low
+ 613.900001n V_low
+ 614.000000n V_low
+ 614.000001n V_hig
+ 614.100000n V_hig
+ 614.100001n V_hig
+ 614.200000n V_hig
+ 614.200001n V_hig
+ 614.300000n V_hig
+ 614.300001n V_hig
+ 614.400000n V_hig
+ 614.400001n V_hig
+ 614.500000n V_hig
+ 614.500001n V_hig
+ 614.600000n V_hig
+ 614.600001n V_hig
+ 614.700000n V_hig
+ 614.700001n V_hig
+ 614.800000n V_hig
+ 614.800001n V_hig
+ 614.900000n V_hig
+ 614.900001n V_hig
+ 615.000000n V_hig
+ 615.000001n V_low
+ 615.100000n V_low
+ 615.100001n V_low
+ 615.200000n V_low
+ 615.200001n V_low
+ 615.300000n V_low
+ 615.300001n V_low
+ 615.400000n V_low
+ 615.400001n V_low
+ 615.500000n V_low
+ 615.500001n V_low
+ 615.600000n V_low
+ 615.600001n V_low
+ 615.700000n V_low
+ 615.700001n V_low
+ 615.800000n V_low
+ 615.800001n V_low
+ 615.900000n V_low
+ 615.900001n V_low
+ 616.000000n V_low
+ 616.000001n V_low
+ 616.100000n V_low
+ 616.100001n V_low
+ 616.200000n V_low
+ 616.200001n V_low
+ 616.300000n V_low
+ 616.300001n V_low
+ 616.400000n V_low
+ 616.400001n V_low
+ 616.500000n V_low
+ 616.500001n V_low
+ 616.600000n V_low
+ 616.600001n V_low
+ 616.700000n V_low
+ 616.700001n V_low
+ 616.800000n V_low
+ 616.800001n V_low
+ 616.900000n V_low
+ 616.900001n V_low
+ 617.000000n V_low
+ 617.000001n V_low
+ 617.100000n V_low
+ 617.100001n V_low
+ 617.200000n V_low
+ 617.200001n V_low
+ 617.300000n V_low
+ 617.300001n V_low
+ 617.400000n V_low
+ 617.400001n V_low
+ 617.500000n V_low
+ 617.500001n V_low
+ 617.600000n V_low
+ 617.600001n V_low
+ 617.700000n V_low
+ 617.700001n V_low
+ 617.800000n V_low
+ 617.800001n V_low
+ 617.900000n V_low
+ 617.900001n V_low
+ 618.000000n V_low
+ 618.000001n V_hig
+ 618.100000n V_hig
+ 618.100001n V_hig
+ 618.200000n V_hig
+ 618.200001n V_hig
+ 618.300000n V_hig
+ 618.300001n V_hig
+ 618.400000n V_hig
+ 618.400001n V_hig
+ 618.500000n V_hig
+ 618.500001n V_hig
+ 618.600000n V_hig
+ 618.600001n V_hig
+ 618.700000n V_hig
+ 618.700001n V_hig
+ 618.800000n V_hig
+ 618.800001n V_hig
+ 618.900000n V_hig
+ 618.900001n V_hig
+ 619.000000n V_hig
+ 619.000001n V_low
+ 619.100000n V_low
+ 619.100001n V_low
+ 619.200000n V_low
+ 619.200001n V_low
+ 619.300000n V_low
+ 619.300001n V_low
+ 619.400000n V_low
+ 619.400001n V_low
+ 619.500000n V_low
+ 619.500001n V_low
+ 619.600000n V_low
+ 619.600001n V_low
+ 619.700000n V_low
+ 619.700001n V_low
+ 619.800000n V_low
+ 619.800001n V_low
+ 619.900000n V_low
+ 619.900001n V_low
+ 620.000000n V_low
+ 620.000001n V_hig
+ 620.100000n V_hig
+ 620.100001n V_hig
+ 620.200000n V_hig
+ 620.200001n V_hig
+ 620.300000n V_hig
+ 620.300001n V_hig
+ 620.400000n V_hig
+ 620.400001n V_hig
+ 620.500000n V_hig
+ 620.500001n V_hig
+ 620.600000n V_hig
+ 620.600001n V_hig
+ 620.700000n V_hig
+ 620.700001n V_hig
+ 620.800000n V_hig
+ 620.800001n V_hig
+ 620.900000n V_hig
+ 620.900001n V_hig
+ 621.000000n V_hig
+ 621.000001n V_hig
+ 621.100000n V_hig
+ 621.100001n V_hig
+ 621.200000n V_hig
+ 621.200001n V_hig
+ 621.300000n V_hig
+ 621.300001n V_hig
+ 621.400000n V_hig
+ 621.400001n V_hig
+ 621.500000n V_hig
+ 621.500001n V_hig
+ 621.600000n V_hig
+ 621.600001n V_hig
+ 621.700000n V_hig
+ 621.700001n V_hig
+ 621.800000n V_hig
+ 621.800001n V_hig
+ 621.900000n V_hig
+ 621.900001n V_hig
+ 622.000000n V_hig
+ 622.000001n V_low
+ 622.100000n V_low
+ 622.100001n V_low
+ 622.200000n V_low
+ 622.200001n V_low
+ 622.300000n V_low
+ 622.300001n V_low
+ 622.400000n V_low
+ 622.400001n V_low
+ 622.500000n V_low
+ 622.500001n V_low
+ 622.600000n V_low
+ 622.600001n V_low
+ 622.700000n V_low
+ 622.700001n V_low
+ 622.800000n V_low
+ 622.800001n V_low
+ 622.900000n V_low
+ 622.900001n V_low
+ 623.000000n V_low
+ 623.000001n V_hig
+ 623.100000n V_hig
+ 623.100001n V_hig
+ 623.200000n V_hig
+ 623.200001n V_hig
+ 623.300000n V_hig
+ 623.300001n V_hig
+ 623.400000n V_hig
+ 623.400001n V_hig
+ 623.500000n V_hig
+ 623.500001n V_hig
+ 623.600000n V_hig
+ 623.600001n V_hig
+ 623.700000n V_hig
+ 623.700001n V_hig
+ 623.800000n V_hig
+ 623.800001n V_hig
+ 623.900000n V_hig
+ 623.900001n V_hig
+ 624.000000n V_hig
+ 624.000001n V_low
+ 624.100000n V_low
+ 624.100001n V_low
+ 624.200000n V_low
+ 624.200001n V_low
+ 624.300000n V_low
+ 624.300001n V_low
+ 624.400000n V_low
+ 624.400001n V_low
+ 624.500000n V_low
+ 624.500001n V_low
+ 624.600000n V_low
+ 624.600001n V_low
+ 624.700000n V_low
+ 624.700001n V_low
+ 624.800000n V_low
+ 624.800001n V_low
+ 624.900000n V_low
+ 624.900001n V_low
+ 625.000000n V_low
+ 625.000001n V_low
+ 625.100000n V_low
+ 625.100001n V_low
+ 625.200000n V_low
+ 625.200001n V_low
+ 625.300000n V_low
+ 625.300001n V_low
+ 625.400000n V_low
+ 625.400001n V_low
+ 625.500000n V_low
+ 625.500001n V_low
+ 625.600000n V_low
+ 625.600001n V_low
+ 625.700000n V_low
+ 625.700001n V_low
+ 625.800000n V_low
+ 625.800001n V_low
+ 625.900000n V_low
+ 625.900001n V_low
+ 626.000000n V_low
+ 626.000001n V_low
+ 626.100000n V_low
+ 626.100001n V_low
+ 626.200000n V_low
+ 626.200001n V_low
+ 626.300000n V_low
+ 626.300001n V_low
+ 626.400000n V_low
+ 626.400001n V_low
+ 626.500000n V_low
+ 626.500001n V_low
+ 626.600000n V_low
+ 626.600001n V_low
+ 626.700000n V_low
+ 626.700001n V_low
+ 626.800000n V_low
+ 626.800001n V_low
+ 626.900000n V_low
+ 626.900001n V_low
+ 627.000000n V_low
+ 627.000001n V_hig
+ 627.100000n V_hig
+ 627.100001n V_hig
+ 627.200000n V_hig
+ 627.200001n V_hig
+ 627.300000n V_hig
+ 627.300001n V_hig
+ 627.400000n V_hig
+ 627.400001n V_hig
+ 627.500000n V_hig
+ 627.500001n V_hig
+ 627.600000n V_hig
+ 627.600001n V_hig
+ 627.700000n V_hig
+ 627.700001n V_hig
+ 627.800000n V_hig
+ 627.800001n V_hig
+ 627.900000n V_hig
+ 627.900001n V_hig
+ 628.000000n V_hig
+ 628.000001n V_low
+ 628.100000n V_low
+ 628.100001n V_low
+ 628.200000n V_low
+ 628.200001n V_low
+ 628.300000n V_low
+ 628.300001n V_low
+ 628.400000n V_low
+ 628.400001n V_low
+ 628.500000n V_low
+ 628.500001n V_low
+ 628.600000n V_low
+ 628.600001n V_low
+ 628.700000n V_low
+ 628.700001n V_low
+ 628.800000n V_low
+ 628.800001n V_low
+ 628.900000n V_low
+ 628.900001n V_low
+ 629.000000n V_low
+ 629.000001n V_low
+ 629.100000n V_low
+ 629.100001n V_low
+ 629.200000n V_low
+ 629.200001n V_low
+ 629.300000n V_low
+ 629.300001n V_low
+ 629.400000n V_low
+ 629.400001n V_low
+ 629.500000n V_low
+ 629.500001n V_low
+ 629.600000n V_low
+ 629.600001n V_low
+ 629.700000n V_low
+ 629.700001n V_low
+ 629.800000n V_low
+ 629.800001n V_low
+ 629.900000n V_low
+ 629.900001n V_low
+ 630.000000n V_low
+ 630.000001n V_low
+ 630.100000n V_low
+ 630.100001n V_low
+ 630.200000n V_low
+ 630.200001n V_low
+ 630.300000n V_low
+ 630.300001n V_low
+ 630.400000n V_low
+ 630.400001n V_low
+ 630.500000n V_low
+ 630.500001n V_low
+ 630.600000n V_low
+ 630.600001n V_low
+ 630.700000n V_low
+ 630.700001n V_low
+ 630.800000n V_low
+ 630.800001n V_low
+ 630.900000n V_low
+ 630.900001n V_low
+ 631.000000n V_low
+ 631.000001n V_hig
+ 631.100000n V_hig
+ 631.100001n V_hig
+ 631.200000n V_hig
+ 631.200001n V_hig
+ 631.300000n V_hig
+ 631.300001n V_hig
+ 631.400000n V_hig
+ 631.400001n V_hig
+ 631.500000n V_hig
+ 631.500001n V_hig
+ 631.600000n V_hig
+ 631.600001n V_hig
+ 631.700000n V_hig
+ 631.700001n V_hig
+ 631.800000n V_hig
+ 631.800001n V_hig
+ 631.900000n V_hig
+ 631.900001n V_hig
+ 632.000000n V_hig
+ 632.000001n V_hig
+ 632.100000n V_hig
+ 632.100001n V_hig
+ 632.200000n V_hig
+ 632.200001n V_hig
+ 632.300000n V_hig
+ 632.300001n V_hig
+ 632.400000n V_hig
+ 632.400001n V_hig
+ 632.500000n V_hig
+ 632.500001n V_hig
+ 632.600000n V_hig
+ 632.600001n V_hig
+ 632.700000n V_hig
+ 632.700001n V_hig
+ 632.800000n V_hig
+ 632.800001n V_hig
+ 632.900000n V_hig
+ 632.900001n V_hig
+ 633.000000n V_hig
+ 633.000001n V_hig
+ 633.100000n V_hig
+ 633.100001n V_hig
+ 633.200000n V_hig
+ 633.200001n V_hig
+ 633.300000n V_hig
+ 633.300001n V_hig
+ 633.400000n V_hig
+ 633.400001n V_hig
+ 633.500000n V_hig
+ 633.500001n V_hig
+ 633.600000n V_hig
+ 633.600001n V_hig
+ 633.700000n V_hig
+ 633.700001n V_hig
+ 633.800000n V_hig
+ 633.800001n V_hig
+ 633.900000n V_hig
+ 633.900001n V_hig
+ 634.000000n V_hig
+ 634.000001n V_hig
+ 634.100000n V_hig
+ 634.100001n V_hig
+ 634.200000n V_hig
+ 634.200001n V_hig
+ 634.300000n V_hig
+ 634.300001n V_hig
+ 634.400000n V_hig
+ 634.400001n V_hig
+ 634.500000n V_hig
+ 634.500001n V_hig
+ 634.600000n V_hig
+ 634.600001n V_hig
+ 634.700000n V_hig
+ 634.700001n V_hig
+ 634.800000n V_hig
+ 634.800001n V_hig
+ 634.900000n V_hig
+ 634.900001n V_hig
+ 635.000000n V_hig
+ 635.000001n V_low
+ 635.100000n V_low
+ 635.100001n V_low
+ 635.200000n V_low
+ 635.200001n V_low
+ 635.300000n V_low
+ 635.300001n V_low
+ 635.400000n V_low
+ 635.400001n V_low
+ 635.500000n V_low
+ 635.500001n V_low
+ 635.600000n V_low
+ 635.600001n V_low
+ 635.700000n V_low
+ 635.700001n V_low
+ 635.800000n V_low
+ 635.800001n V_low
+ 635.900000n V_low
+ 635.900001n V_low
+ 636.000000n V_low
+ 636.000001n V_hig
+ 636.100000n V_hig
+ 636.100001n V_hig
+ 636.200000n V_hig
+ 636.200001n V_hig
+ 636.300000n V_hig
+ 636.300001n V_hig
+ 636.400000n V_hig
+ 636.400001n V_hig
+ 636.500000n V_hig
+ 636.500001n V_hig
+ 636.600000n V_hig
+ 636.600001n V_hig
+ 636.700000n V_hig
+ 636.700001n V_hig
+ 636.800000n V_hig
+ 636.800001n V_hig
+ 636.900000n V_hig
+ 636.900001n V_hig
+ 637.000000n V_hig
+ 637.000001n V_hig
+ 637.100000n V_hig
+ 637.100001n V_hig
+ 637.200000n V_hig
+ 637.200001n V_hig
+ 637.300000n V_hig
+ 637.300001n V_hig
+ 637.400000n V_hig
+ 637.400001n V_hig
+ 637.500000n V_hig
+ 637.500001n V_hig
+ 637.600000n V_hig
+ 637.600001n V_hig
+ 637.700000n V_hig
+ 637.700001n V_hig
+ 637.800000n V_hig
+ 637.800001n V_hig
+ 637.900000n V_hig
+ 637.900001n V_hig
+ 638.000000n V_hig
+ 638.000001n V_low
+ 638.100000n V_low
+ 638.100001n V_low
+ 638.200000n V_low
+ 638.200001n V_low
+ 638.300000n V_low
+ 638.300001n V_low
+ 638.400000n V_low
+ 638.400001n V_low
+ 638.500000n V_low
+ 638.500001n V_low
+ 638.600000n V_low
+ 638.600001n V_low
+ 638.700000n V_low
+ 638.700001n V_low
+ 638.800000n V_low
+ 638.800001n V_low
+ 638.900000n V_low
+ 638.900001n V_low
+ 639.000000n V_low
+ 639.000001n V_low
+ 639.100000n V_low
+ 639.100001n V_low
+ 639.200000n V_low
+ 639.200001n V_low
+ 639.300000n V_low
+ 639.300001n V_low
+ 639.400000n V_low
+ 639.400001n V_low
+ 639.500000n V_low
+ 639.500001n V_low
+ 639.600000n V_low
+ 639.600001n V_low
+ 639.700000n V_low
+ 639.700001n V_low
+ 639.800000n V_low
+ 639.800001n V_low
+ 639.900000n V_low
+ 639.900001n V_low
+ 640.000000n V_low
+ 640.000001n V_hig
+ 640.100000n V_hig
+ 640.100001n V_hig
+ 640.200000n V_hig
+ 640.200001n V_hig
+ 640.300000n V_hig
+ 640.300001n V_hig
+ 640.400000n V_hig
+ 640.400001n V_hig
+ 640.500000n V_hig
+ 640.500001n V_hig
+ 640.600000n V_hig
+ 640.600001n V_hig
+ 640.700000n V_hig
+ 640.700001n V_hig
+ 640.800000n V_hig
+ 640.800001n V_hig
+ 640.900000n V_hig
+ 640.900001n V_hig
+ 641.000000n V_hig
+ 641.000001n V_hig
+ 641.100000n V_hig
+ 641.100001n V_hig
+ 641.200000n V_hig
+ 641.200001n V_hig
+ 641.300000n V_hig
+ 641.300001n V_hig
+ 641.400000n V_hig
+ 641.400001n V_hig
+ 641.500000n V_hig
+ 641.500001n V_hig
+ 641.600000n V_hig
+ 641.600001n V_hig
+ 641.700000n V_hig
+ 641.700001n V_hig
+ 641.800000n V_hig
+ 641.800001n V_hig
+ 641.900000n V_hig
+ 641.900001n V_hig
+ 642.000000n V_hig
+ 642.000001n V_low
+ 642.100000n V_low
+ 642.100001n V_low
+ 642.200000n V_low
+ 642.200001n V_low
+ 642.300000n V_low
+ 642.300001n V_low
+ 642.400000n V_low
+ 642.400001n V_low
+ 642.500000n V_low
+ 642.500001n V_low
+ 642.600000n V_low
+ 642.600001n V_low
+ 642.700000n V_low
+ 642.700001n V_low
+ 642.800000n V_low
+ 642.800001n V_low
+ 642.900000n V_low
+ 642.900001n V_low
+ 643.000000n V_low
+ 643.000001n V_hig
+ 643.100000n V_hig
+ 643.100001n V_hig
+ 643.200000n V_hig
+ 643.200001n V_hig
+ 643.300000n V_hig
+ 643.300001n V_hig
+ 643.400000n V_hig
+ 643.400001n V_hig
+ 643.500000n V_hig
+ 643.500001n V_hig
+ 643.600000n V_hig
+ 643.600001n V_hig
+ 643.700000n V_hig
+ 643.700001n V_hig
+ 643.800000n V_hig
+ 643.800001n V_hig
+ 643.900000n V_hig
+ 643.900001n V_hig
+ 644.000000n V_hig
+ 644.000001n V_low
+ 644.100000n V_low
+ 644.100001n V_low
+ 644.200000n V_low
+ 644.200001n V_low
+ 644.300000n V_low
+ 644.300001n V_low
+ 644.400000n V_low
+ 644.400001n V_low
+ 644.500000n V_low
+ 644.500001n V_low
+ 644.600000n V_low
+ 644.600001n V_low
+ 644.700000n V_low
+ 644.700001n V_low
+ 644.800000n V_low
+ 644.800001n V_low
+ 644.900000n V_low
+ 644.900001n V_low
+ 645.000000n V_low
+ 645.000001n V_low
+ 645.100000n V_low
+ 645.100001n V_low
+ 645.200000n V_low
+ 645.200001n V_low
+ 645.300000n V_low
+ 645.300001n V_low
+ 645.400000n V_low
+ 645.400001n V_low
+ 645.500000n V_low
+ 645.500001n V_low
+ 645.600000n V_low
+ 645.600001n V_low
+ 645.700000n V_low
+ 645.700001n V_low
+ 645.800000n V_low
+ 645.800001n V_low
+ 645.900000n V_low
+ 645.900001n V_low
+ 646.000000n V_low
+ 646.000001n V_hig
+ 646.100000n V_hig
+ 646.100001n V_hig
+ 646.200000n V_hig
+ 646.200001n V_hig
+ 646.300000n V_hig
+ 646.300001n V_hig
+ 646.400000n V_hig
+ 646.400001n V_hig
+ 646.500000n V_hig
+ 646.500001n V_hig
+ 646.600000n V_hig
+ 646.600001n V_hig
+ 646.700000n V_hig
+ 646.700001n V_hig
+ 646.800000n V_hig
+ 646.800001n V_hig
+ 646.900000n V_hig
+ 646.900001n V_hig
+ 647.000000n V_hig
+ 647.000001n V_low
+ 647.100000n V_low
+ 647.100001n V_low
+ 647.200000n V_low
+ 647.200001n V_low
+ 647.300000n V_low
+ 647.300001n V_low
+ 647.400000n V_low
+ 647.400001n V_low
+ 647.500000n V_low
+ 647.500001n V_low
+ 647.600000n V_low
+ 647.600001n V_low
+ 647.700000n V_low
+ 647.700001n V_low
+ 647.800000n V_low
+ 647.800001n V_low
+ 647.900000n V_low
+ 647.900001n V_low
+ 648.000000n V_low
+ 648.000001n V_hig
+ 648.100000n V_hig
+ 648.100001n V_hig
+ 648.200000n V_hig
+ 648.200001n V_hig
+ 648.300000n V_hig
+ 648.300001n V_hig
+ 648.400000n V_hig
+ 648.400001n V_hig
+ 648.500000n V_hig
+ 648.500001n V_hig
+ 648.600000n V_hig
+ 648.600001n V_hig
+ 648.700000n V_hig
+ 648.700001n V_hig
+ 648.800000n V_hig
+ 648.800001n V_hig
+ 648.900000n V_hig
+ 648.900001n V_hig
+ 649.000000n V_hig
+ 649.000001n V_hig
+ 649.100000n V_hig
+ 649.100001n V_hig
+ 649.200000n V_hig
+ 649.200001n V_hig
+ 649.300000n V_hig
+ 649.300001n V_hig
+ 649.400000n V_hig
+ 649.400001n V_hig
+ 649.500000n V_hig
+ 649.500001n V_hig
+ 649.600000n V_hig
+ 649.600001n V_hig
+ 649.700000n V_hig
+ 649.700001n V_hig
+ 649.800000n V_hig
+ 649.800001n V_hig
+ 649.900000n V_hig
+ 649.900001n V_hig
+ 650.000000n V_hig
+ 650.000001n V_hig
+ 650.100000n V_hig
+ 650.100001n V_hig
+ 650.200000n V_hig
+ 650.200001n V_hig
+ 650.300000n V_hig
+ 650.300001n V_hig
+ 650.400000n V_hig
+ 650.400001n V_hig
+ 650.500000n V_hig
+ 650.500001n V_hig
+ 650.600000n V_hig
+ 650.600001n V_hig
+ 650.700000n V_hig
+ 650.700001n V_hig
+ 650.800000n V_hig
+ 650.800001n V_hig
+ 650.900000n V_hig
+ 650.900001n V_hig
+ 651.000000n V_hig
+ 651.000001n V_hig
+ 651.100000n V_hig
+ 651.100001n V_hig
+ 651.200000n V_hig
+ 651.200001n V_hig
+ 651.300000n V_hig
+ 651.300001n V_hig
+ 651.400000n V_hig
+ 651.400001n V_hig
+ 651.500000n V_hig
+ 651.500001n V_hig
+ 651.600000n V_hig
+ 651.600001n V_hig
+ 651.700000n V_hig
+ 651.700001n V_hig
+ 651.800000n V_hig
+ 651.800001n V_hig
+ 651.900000n V_hig
+ 651.900001n V_hig
+ 652.000000n V_hig
+ 652.000001n V_hig
+ 652.100000n V_hig
+ 652.100001n V_hig
+ 652.200000n V_hig
+ 652.200001n V_hig
+ 652.300000n V_hig
+ 652.300001n V_hig
+ 652.400000n V_hig
+ 652.400001n V_hig
+ 652.500000n V_hig
+ 652.500001n V_hig
+ 652.600000n V_hig
+ 652.600001n V_hig
+ 652.700000n V_hig
+ 652.700001n V_hig
+ 652.800000n V_hig
+ 652.800001n V_hig
+ 652.900000n V_hig
+ 652.900001n V_hig
+ 653.000000n V_hig
+ 653.000001n V_low
+ 653.100000n V_low
+ 653.100001n V_low
+ 653.200000n V_low
+ 653.200001n V_low
+ 653.300000n V_low
+ 653.300001n V_low
+ 653.400000n V_low
+ 653.400001n V_low
+ 653.500000n V_low
+ 653.500001n V_low
+ 653.600000n V_low
+ 653.600001n V_low
+ 653.700000n V_low
+ 653.700001n V_low
+ 653.800000n V_low
+ 653.800001n V_low
+ 653.900000n V_low
+ 653.900001n V_low
+ 654.000000n V_low
+ 654.000001n V_hig
+ 654.100000n V_hig
+ 654.100001n V_hig
+ 654.200000n V_hig
+ 654.200001n V_hig
+ 654.300000n V_hig
+ 654.300001n V_hig
+ 654.400000n V_hig
+ 654.400001n V_hig
+ 654.500000n V_hig
+ 654.500001n V_hig
+ 654.600000n V_hig
+ 654.600001n V_hig
+ 654.700000n V_hig
+ 654.700001n V_hig
+ 654.800000n V_hig
+ 654.800001n V_hig
+ 654.900000n V_hig
+ 654.900001n V_hig
+ 655.000000n V_hig
+ 655.000001n V_hig
+ 655.100000n V_hig
+ 655.100001n V_hig
+ 655.200000n V_hig
+ 655.200001n V_hig
+ 655.300000n V_hig
+ 655.300001n V_hig
+ 655.400000n V_hig
+ 655.400001n V_hig
+ 655.500000n V_hig
+ 655.500001n V_hig
+ 655.600000n V_hig
+ 655.600001n V_hig
+ 655.700000n V_hig
+ 655.700001n V_hig
+ 655.800000n V_hig
+ 655.800001n V_hig
+ 655.900000n V_hig
+ 655.900001n V_hig
+ 656.000000n V_hig
+ 656.000001n V_low
+ 656.100000n V_low
+ 656.100001n V_low
+ 656.200000n V_low
+ 656.200001n V_low
+ 656.300000n V_low
+ 656.300001n V_low
+ 656.400000n V_low
+ 656.400001n V_low
+ 656.500000n V_low
+ 656.500001n V_low
+ 656.600000n V_low
+ 656.600001n V_low
+ 656.700000n V_low
+ 656.700001n V_low
+ 656.800000n V_low
+ 656.800001n V_low
+ 656.900000n V_low
+ 656.900001n V_low
+ 657.000000n V_low
+ 657.000001n V_low
+ 657.100000n V_low
+ 657.100001n V_low
+ 657.200000n V_low
+ 657.200001n V_low
+ 657.300000n V_low
+ 657.300001n V_low
+ 657.400000n V_low
+ 657.400001n V_low
+ 657.500000n V_low
+ 657.500001n V_low
+ 657.600000n V_low
+ 657.600001n V_low
+ 657.700000n V_low
+ 657.700001n V_low
+ 657.800000n V_low
+ 657.800001n V_low
+ 657.900000n V_low
+ 657.900001n V_low
+ 658.000000n V_low
+ 658.000001n V_hig
+ 658.100000n V_hig
+ 658.100001n V_hig
+ 658.200000n V_hig
+ 658.200001n V_hig
+ 658.300000n V_hig
+ 658.300001n V_hig
+ 658.400000n V_hig
+ 658.400001n V_hig
+ 658.500000n V_hig
+ 658.500001n V_hig
+ 658.600000n V_hig
+ 658.600001n V_hig
+ 658.700000n V_hig
+ 658.700001n V_hig
+ 658.800000n V_hig
+ 658.800001n V_hig
+ 658.900000n V_hig
+ 658.900001n V_hig
+ 659.000000n V_hig
+ 659.000001n V_hig
+ 659.100000n V_hig
+ 659.100001n V_hig
+ 659.200000n V_hig
+ 659.200001n V_hig
+ 659.300000n V_hig
+ 659.300001n V_hig
+ 659.400000n V_hig
+ 659.400001n V_hig
+ 659.500000n V_hig
+ 659.500001n V_hig
+ 659.600000n V_hig
+ 659.600001n V_hig
+ 659.700000n V_hig
+ 659.700001n V_hig
+ 659.800000n V_hig
+ 659.800001n V_hig
+ 659.900000n V_hig
+ 659.900001n V_hig
+ 660.000000n V_hig
+ 660.000001n V_low
+ 660.100000n V_low
+ 660.100001n V_low
+ 660.200000n V_low
+ 660.200001n V_low
+ 660.300000n V_low
+ 660.300001n V_low
+ 660.400000n V_low
+ 660.400001n V_low
+ 660.500000n V_low
+ 660.500001n V_low
+ 660.600000n V_low
+ 660.600001n V_low
+ 660.700000n V_low
+ 660.700001n V_low
+ 660.800000n V_low
+ 660.800001n V_low
+ 660.900000n V_low
+ 660.900001n V_low
+ 661.000000n V_low
+ 661.000001n V_low
+ 661.100000n V_low
+ 661.100001n V_low
+ 661.200000n V_low
+ 661.200001n V_low
+ 661.300000n V_low
+ 661.300001n V_low
+ 661.400000n V_low
+ 661.400001n V_low
+ 661.500000n V_low
+ 661.500001n V_low
+ 661.600000n V_low
+ 661.600001n V_low
+ 661.700000n V_low
+ 661.700001n V_low
+ 661.800000n V_low
+ 661.800001n V_low
+ 661.900000n V_low
+ 661.900001n V_low
+ 662.000000n V_low
+ 662.000001n V_low
+ 662.100000n V_low
+ 662.100001n V_low
+ 662.200000n V_low
+ 662.200001n V_low
+ 662.300000n V_low
+ 662.300001n V_low
+ 662.400000n V_low
+ 662.400001n V_low
+ 662.500000n V_low
+ 662.500001n V_low
+ 662.600000n V_low
+ 662.600001n V_low
+ 662.700000n V_low
+ 662.700001n V_low
+ 662.800000n V_low
+ 662.800001n V_low
+ 662.900000n V_low
+ 662.900001n V_low
+ 663.000000n V_low
+ 663.000001n V_low
+ 663.100000n V_low
+ 663.100001n V_low
+ 663.200000n V_low
+ 663.200001n V_low
+ 663.300000n V_low
+ 663.300001n V_low
+ 663.400000n V_low
+ 663.400001n V_low
+ 663.500000n V_low
+ 663.500001n V_low
+ 663.600000n V_low
+ 663.600001n V_low
+ 663.700000n V_low
+ 663.700001n V_low
+ 663.800000n V_low
+ 663.800001n V_low
+ 663.900000n V_low
+ 663.900001n V_low
+ 664.000000n V_low
+ 664.000001n V_low
+ 664.100000n V_low
+ 664.100001n V_low
+ 664.200000n V_low
+ 664.200001n V_low
+ 664.300000n V_low
+ 664.300001n V_low
+ 664.400000n V_low
+ 664.400001n V_low
+ 664.500000n V_low
+ 664.500001n V_low
+ 664.600000n V_low
+ 664.600001n V_low
+ 664.700000n V_low
+ 664.700001n V_low
+ 664.800000n V_low
+ 664.800001n V_low
+ 664.900000n V_low
+ 664.900001n V_low
+ 665.000000n V_low
+ 665.000001n V_hig
+ 665.100000n V_hig
+ 665.100001n V_hig
+ 665.200000n V_hig
+ 665.200001n V_hig
+ 665.300000n V_hig
+ 665.300001n V_hig
+ 665.400000n V_hig
+ 665.400001n V_hig
+ 665.500000n V_hig
+ 665.500001n V_hig
+ 665.600000n V_hig
+ 665.600001n V_hig
+ 665.700000n V_hig
+ 665.700001n V_hig
+ 665.800000n V_hig
+ 665.800001n V_hig
+ 665.900000n V_hig
+ 665.900001n V_hig
+ 666.000000n V_hig
+ 666.000001n V_low
+ 666.100000n V_low
+ 666.100001n V_low
+ 666.200000n V_low
+ 666.200001n V_low
+ 666.300000n V_low
+ 666.300001n V_low
+ 666.400000n V_low
+ 666.400001n V_low
+ 666.500000n V_low
+ 666.500001n V_low
+ 666.600000n V_low
+ 666.600001n V_low
+ 666.700000n V_low
+ 666.700001n V_low
+ 666.800000n V_low
+ 666.800001n V_low
+ 666.900000n V_low
+ 666.900001n V_low
+ 667.000000n V_low
+ 667.000001n V_low
+ 667.100000n V_low
+ 667.100001n V_low
+ 667.200000n V_low
+ 667.200001n V_low
+ 667.300000n V_low
+ 667.300001n V_low
+ 667.400000n V_low
+ 667.400001n V_low
+ 667.500000n V_low
+ 667.500001n V_low
+ 667.600000n V_low
+ 667.600001n V_low
+ 667.700000n V_low
+ 667.700001n V_low
+ 667.800000n V_low
+ 667.800001n V_low
+ 667.900000n V_low
+ 667.900001n V_low
+ 668.000000n V_low
+ 668.000001n V_low
+ 668.100000n V_low
+ 668.100001n V_low
+ 668.200000n V_low
+ 668.200001n V_low
+ 668.300000n V_low
+ 668.300001n V_low
+ 668.400000n V_low
+ 668.400001n V_low
+ 668.500000n V_low
+ 668.500001n V_low
+ 668.600000n V_low
+ 668.600001n V_low
+ 668.700000n V_low
+ 668.700001n V_low
+ 668.800000n V_low
+ 668.800001n V_low
+ 668.900000n V_low
+ 668.900001n V_low
+ 669.000000n V_low
+ 669.000001n V_low
+ 669.100000n V_low
+ 669.100001n V_low
+ 669.200000n V_low
+ 669.200001n V_low
+ 669.300000n V_low
+ 669.300001n V_low
+ 669.400000n V_low
+ 669.400001n V_low
+ 669.500000n V_low
+ 669.500001n V_low
+ 669.600000n V_low
+ 669.600001n V_low
+ 669.700000n V_low
+ 669.700001n V_low
+ 669.800000n V_low
+ 669.800001n V_low
+ 669.900000n V_low
+ 669.900001n V_low
+ 670.000000n V_low
+ 670.000001n V_hig
+ 670.100000n V_hig
+ 670.100001n V_hig
+ 670.200000n V_hig
+ 670.200001n V_hig
+ 670.300000n V_hig
+ 670.300001n V_hig
+ 670.400000n V_hig
+ 670.400001n V_hig
+ 670.500000n V_hig
+ 670.500001n V_hig
+ 670.600000n V_hig
+ 670.600001n V_hig
+ 670.700000n V_hig
+ 670.700001n V_hig
+ 670.800000n V_hig
+ 670.800001n V_hig
+ 670.900000n V_hig
+ 670.900001n V_hig
+ 671.000000n V_hig
+ 671.000001n V_hig
+ 671.100000n V_hig
+ 671.100001n V_hig
+ 671.200000n V_hig
+ 671.200001n V_hig
+ 671.300000n V_hig
+ 671.300001n V_hig
+ 671.400000n V_hig
+ 671.400001n V_hig
+ 671.500000n V_hig
+ 671.500001n V_hig
+ 671.600000n V_hig
+ 671.600001n V_hig
+ 671.700000n V_hig
+ 671.700001n V_hig
+ 671.800000n V_hig
+ 671.800001n V_hig
+ 671.900000n V_hig
+ 671.900001n V_hig
+ 672.000000n V_hig
+ 672.000001n V_hig
+ 672.100000n V_hig
+ 672.100001n V_hig
+ 672.200000n V_hig
+ 672.200001n V_hig
+ 672.300000n V_hig
+ 672.300001n V_hig
+ 672.400000n V_hig
+ 672.400001n V_hig
+ 672.500000n V_hig
+ 672.500001n V_hig
+ 672.600000n V_hig
+ 672.600001n V_hig
+ 672.700000n V_hig
+ 672.700001n V_hig
+ 672.800000n V_hig
+ 672.800001n V_hig
+ 672.900000n V_hig
+ 672.900001n V_hig
+ 673.000000n V_hig
+ 673.000001n V_low
+ 673.100000n V_low
+ 673.100001n V_low
+ 673.200000n V_low
+ 673.200001n V_low
+ 673.300000n V_low
+ 673.300001n V_low
+ 673.400000n V_low
+ 673.400001n V_low
+ 673.500000n V_low
+ 673.500001n V_low
+ 673.600000n V_low
+ 673.600001n V_low
+ 673.700000n V_low
+ 673.700001n V_low
+ 673.800000n V_low
+ 673.800001n V_low
+ 673.900000n V_low
+ 673.900001n V_low
+ 674.000000n V_low
+ 674.000001n V_hig
+ 674.100000n V_hig
+ 674.100001n V_hig
+ 674.200000n V_hig
+ 674.200001n V_hig
+ 674.300000n V_hig
+ 674.300001n V_hig
+ 674.400000n V_hig
+ 674.400001n V_hig
+ 674.500000n V_hig
+ 674.500001n V_hig
+ 674.600000n V_hig
+ 674.600001n V_hig
+ 674.700000n V_hig
+ 674.700001n V_hig
+ 674.800000n V_hig
+ 674.800001n V_hig
+ 674.900000n V_hig
+ 674.900001n V_hig
+ 675.000000n V_hig
+ 675.000001n V_hig
+ 675.100000n V_hig
+ 675.100001n V_hig
+ 675.200000n V_hig
+ 675.200001n V_hig
+ 675.300000n V_hig
+ 675.300001n V_hig
+ 675.400000n V_hig
+ 675.400001n V_hig
+ 675.500000n V_hig
+ 675.500001n V_hig
+ 675.600000n V_hig
+ 675.600001n V_hig
+ 675.700000n V_hig
+ 675.700001n V_hig
+ 675.800000n V_hig
+ 675.800001n V_hig
+ 675.900000n V_hig
+ 675.900001n V_hig
+ 676.000000n V_hig
+ 676.000001n V_low
+ 676.100000n V_low
+ 676.100001n V_low
+ 676.200000n V_low
+ 676.200001n V_low
+ 676.300000n V_low
+ 676.300001n V_low
+ 676.400000n V_low
+ 676.400001n V_low
+ 676.500000n V_low
+ 676.500001n V_low
+ 676.600000n V_low
+ 676.600001n V_low
+ 676.700000n V_low
+ 676.700001n V_low
+ 676.800000n V_low
+ 676.800001n V_low
+ 676.900000n V_low
+ 676.900001n V_low
+ 677.000000n V_low
+ 677.000001n V_hig
+ 677.100000n V_hig
+ 677.100001n V_hig
+ 677.200000n V_hig
+ 677.200001n V_hig
+ 677.300000n V_hig
+ 677.300001n V_hig
+ 677.400000n V_hig
+ 677.400001n V_hig
+ 677.500000n V_hig
+ 677.500001n V_hig
+ 677.600000n V_hig
+ 677.600001n V_hig
+ 677.700000n V_hig
+ 677.700001n V_hig
+ 677.800000n V_hig
+ 677.800001n V_hig
+ 677.900000n V_hig
+ 677.900001n V_hig
+ 678.000000n V_hig
+ 678.000001n V_hig
+ 678.100000n V_hig
+ 678.100001n V_hig
+ 678.200000n V_hig
+ 678.200001n V_hig
+ 678.300000n V_hig
+ 678.300001n V_hig
+ 678.400000n V_hig
+ 678.400001n V_hig
+ 678.500000n V_hig
+ 678.500001n V_hig
+ 678.600000n V_hig
+ 678.600001n V_hig
+ 678.700000n V_hig
+ 678.700001n V_hig
+ 678.800000n V_hig
+ 678.800001n V_hig
+ 678.900000n V_hig
+ 678.900001n V_hig
+ 679.000000n V_hig
+ 679.000001n V_hig
+ 679.100000n V_hig
+ 679.100001n V_hig
+ 679.200000n V_hig
+ 679.200001n V_hig
+ 679.300000n V_hig
+ 679.300001n V_hig
+ 679.400000n V_hig
+ 679.400001n V_hig
+ 679.500000n V_hig
+ 679.500001n V_hig
+ 679.600000n V_hig
+ 679.600001n V_hig
+ 679.700000n V_hig
+ 679.700001n V_hig
+ 679.800000n V_hig
+ 679.800001n V_hig
+ 679.900000n V_hig
+ 679.900001n V_hig
+ 680.000000n V_hig
+ 680.000001n V_hig
+ 680.100000n V_hig
+ 680.100001n V_hig
+ 680.200000n V_hig
+ 680.200001n V_hig
+ 680.300000n V_hig
+ 680.300001n V_hig
+ 680.400000n V_hig
+ 680.400001n V_hig
+ 680.500000n V_hig
+ 680.500001n V_hig
+ 680.600000n V_hig
+ 680.600001n V_hig
+ 680.700000n V_hig
+ 680.700001n V_hig
+ 680.800000n V_hig
+ 680.800001n V_hig
+ 680.900000n V_hig
+ 680.900001n V_hig
+ 681.000000n V_hig
+ 681.000001n V_hig
+ 681.100000n V_hig
+ 681.100001n V_hig
+ 681.200000n V_hig
+ 681.200001n V_hig
+ 681.300000n V_hig
+ 681.300001n V_hig
+ 681.400000n V_hig
+ 681.400001n V_hig
+ 681.500000n V_hig
+ 681.500001n V_hig
+ 681.600000n V_hig
+ 681.600001n V_hig
+ 681.700000n V_hig
+ 681.700001n V_hig
+ 681.800000n V_hig
+ 681.800001n V_hig
+ 681.900000n V_hig
+ 681.900001n V_hig
+ 682.000000n V_hig
+ 682.000001n V_hig
+ 682.100000n V_hig
+ 682.100001n V_hig
+ 682.200000n V_hig
+ 682.200001n V_hig
+ 682.300000n V_hig
+ 682.300001n V_hig
+ 682.400000n V_hig
+ 682.400001n V_hig
+ 682.500000n V_hig
+ 682.500001n V_hig
+ 682.600000n V_hig
+ 682.600001n V_hig
+ 682.700000n V_hig
+ 682.700001n V_hig
+ 682.800000n V_hig
+ 682.800001n V_hig
+ 682.900000n V_hig
+ 682.900001n V_hig
+ 683.000000n V_hig
+ 683.000001n V_low
+ 683.100000n V_low
+ 683.100001n V_low
+ 683.200000n V_low
+ 683.200001n V_low
+ 683.300000n V_low
+ 683.300001n V_low
+ 683.400000n V_low
+ 683.400001n V_low
+ 683.500000n V_low
+ 683.500001n V_low
+ 683.600000n V_low
+ 683.600001n V_low
+ 683.700000n V_low
+ 683.700001n V_low
+ 683.800000n V_low
+ 683.800001n V_low
+ 683.900000n V_low
+ 683.900001n V_low
+ 684.000000n V_low
+ 684.000001n V_hig
+ 684.100000n V_hig
+ 684.100001n V_hig
+ 684.200000n V_hig
+ 684.200001n V_hig
+ 684.300000n V_hig
+ 684.300001n V_hig
+ 684.400000n V_hig
+ 684.400001n V_hig
+ 684.500000n V_hig
+ 684.500001n V_hig
+ 684.600000n V_hig
+ 684.600001n V_hig
+ 684.700000n V_hig
+ 684.700001n V_hig
+ 684.800000n V_hig
+ 684.800001n V_hig
+ 684.900000n V_hig
+ 684.900001n V_hig
+ 685.000000n V_hig
+ 685.000001n V_low
+ 685.100000n V_low
+ 685.100001n V_low
+ 685.200000n V_low
+ 685.200001n V_low
+ 685.300000n V_low
+ 685.300001n V_low
+ 685.400000n V_low
+ 685.400001n V_low
+ 685.500000n V_low
+ 685.500001n V_low
+ 685.600000n V_low
+ 685.600001n V_low
+ 685.700000n V_low
+ 685.700001n V_low
+ 685.800000n V_low
+ 685.800001n V_low
+ 685.900000n V_low
+ 685.900001n V_low
+ 686.000000n V_low
+ 686.000001n V_hig
+ 686.100000n V_hig
+ 686.100001n V_hig
+ 686.200000n V_hig
+ 686.200001n V_hig
+ 686.300000n V_hig
+ 686.300001n V_hig
+ 686.400000n V_hig
+ 686.400001n V_hig
+ 686.500000n V_hig
+ 686.500001n V_hig
+ 686.600000n V_hig
+ 686.600001n V_hig
+ 686.700000n V_hig
+ 686.700001n V_hig
+ 686.800000n V_hig
+ 686.800001n V_hig
+ 686.900000n V_hig
+ 686.900001n V_hig
+ 687.000000n V_hig
+ 687.000001n V_low
+ 687.100000n V_low
+ 687.100001n V_low
+ 687.200000n V_low
+ 687.200001n V_low
+ 687.300000n V_low
+ 687.300001n V_low
+ 687.400000n V_low
+ 687.400001n V_low
+ 687.500000n V_low
+ 687.500001n V_low
+ 687.600000n V_low
+ 687.600001n V_low
+ 687.700000n V_low
+ 687.700001n V_low
+ 687.800000n V_low
+ 687.800001n V_low
+ 687.900000n V_low
+ 687.900001n V_low
+ 688.000000n V_low
+ 688.000001n V_hig
+ 688.100000n V_hig
+ 688.100001n V_hig
+ 688.200000n V_hig
+ 688.200001n V_hig
+ 688.300000n V_hig
+ 688.300001n V_hig
+ 688.400000n V_hig
+ 688.400001n V_hig
+ 688.500000n V_hig
+ 688.500001n V_hig
+ 688.600000n V_hig
+ 688.600001n V_hig
+ 688.700000n V_hig
+ 688.700001n V_hig
+ 688.800000n V_hig
+ 688.800001n V_hig
+ 688.900000n V_hig
+ 688.900001n V_hig
+ 689.000000n V_hig
+ 689.000001n V_low
+ 689.100000n V_low
+ 689.100001n V_low
+ 689.200000n V_low
+ 689.200001n V_low
+ 689.300000n V_low
+ 689.300001n V_low
+ 689.400000n V_low
+ 689.400001n V_low
+ 689.500000n V_low
+ 689.500001n V_low
+ 689.600000n V_low
+ 689.600001n V_low
+ 689.700000n V_low
+ 689.700001n V_low
+ 689.800000n V_low
+ 689.800001n V_low
+ 689.900000n V_low
+ 689.900001n V_low
+ 690.000000n V_low
+ 690.000001n V_hig
+ 690.100000n V_hig
+ 690.100001n V_hig
+ 690.200000n V_hig
+ 690.200001n V_hig
+ 690.300000n V_hig
+ 690.300001n V_hig
+ 690.400000n V_hig
+ 690.400001n V_hig
+ 690.500000n V_hig
+ 690.500001n V_hig
+ 690.600000n V_hig
+ 690.600001n V_hig
+ 690.700000n V_hig
+ 690.700001n V_hig
+ 690.800000n V_hig
+ 690.800001n V_hig
+ 690.900000n V_hig
+ 690.900001n V_hig
+ 691.000000n V_hig
+ 691.000001n V_hig
+ 691.100000n V_hig
+ 691.100001n V_hig
+ 691.200000n V_hig
+ 691.200001n V_hig
+ 691.300000n V_hig
+ 691.300001n V_hig
+ 691.400000n V_hig
+ 691.400001n V_hig
+ 691.500000n V_hig
+ 691.500001n V_hig
+ 691.600000n V_hig
+ 691.600001n V_hig
+ 691.700000n V_hig
+ 691.700001n V_hig
+ 691.800000n V_hig
+ 691.800001n V_hig
+ 691.900000n V_hig
+ 691.900001n V_hig
+ 692.000000n V_hig
+ 692.000001n V_low
+ 692.100000n V_low
+ 692.100001n V_low
+ 692.200000n V_low
+ 692.200001n V_low
+ 692.300000n V_low
+ 692.300001n V_low
+ 692.400000n V_low
+ 692.400001n V_low
+ 692.500000n V_low
+ 692.500001n V_low
+ 692.600000n V_low
+ 692.600001n V_low
+ 692.700000n V_low
+ 692.700001n V_low
+ 692.800000n V_low
+ 692.800001n V_low
+ 692.900000n V_low
+ 692.900001n V_low
+ 693.000000n V_low
+ 693.000001n V_hig
+ 693.100000n V_hig
+ 693.100001n V_hig
+ 693.200000n V_hig
+ 693.200001n V_hig
+ 693.300000n V_hig
+ 693.300001n V_hig
+ 693.400000n V_hig
+ 693.400001n V_hig
+ 693.500000n V_hig
+ 693.500001n V_hig
+ 693.600000n V_hig
+ 693.600001n V_hig
+ 693.700000n V_hig
+ 693.700001n V_hig
+ 693.800000n V_hig
+ 693.800001n V_hig
+ 693.900000n V_hig
+ 693.900001n V_hig
+ 694.000000n V_hig
+ 694.000001n V_hig
+ 694.100000n V_hig
+ 694.100001n V_hig
+ 694.200000n V_hig
+ 694.200001n V_hig
+ 694.300000n V_hig
+ 694.300001n V_hig
+ 694.400000n V_hig
+ 694.400001n V_hig
+ 694.500000n V_hig
+ 694.500001n V_hig
+ 694.600000n V_hig
+ 694.600001n V_hig
+ 694.700000n V_hig
+ 694.700001n V_hig
+ 694.800000n V_hig
+ 694.800001n V_hig
+ 694.900000n V_hig
+ 694.900001n V_hig
+ 695.000000n V_hig
+ 695.000001n V_hig
+ 695.100000n V_hig
+ 695.100001n V_hig
+ 695.200000n V_hig
+ 695.200001n V_hig
+ 695.300000n V_hig
+ 695.300001n V_hig
+ 695.400000n V_hig
+ 695.400001n V_hig
+ 695.500000n V_hig
+ 695.500001n V_hig
+ 695.600000n V_hig
+ 695.600001n V_hig
+ 695.700000n V_hig
+ 695.700001n V_hig
+ 695.800000n V_hig
+ 695.800001n V_hig
+ 695.900000n V_hig
+ 695.900001n V_hig
+ 696.000000n V_hig
+ 696.000001n V_low
+ 696.100000n V_low
+ 696.100001n V_low
+ 696.200000n V_low
+ 696.200001n V_low
+ 696.300000n V_low
+ 696.300001n V_low
+ 696.400000n V_low
+ 696.400001n V_low
+ 696.500000n V_low
+ 696.500001n V_low
+ 696.600000n V_low
+ 696.600001n V_low
+ 696.700000n V_low
+ 696.700001n V_low
+ 696.800000n V_low
+ 696.800001n V_low
+ 696.900000n V_low
+ 696.900001n V_low
+ 697.000000n V_low
+ 697.000001n V_hig
+ 697.100000n V_hig
+ 697.100001n V_hig
+ 697.200000n V_hig
+ 697.200001n V_hig
+ 697.300000n V_hig
+ 697.300001n V_hig
+ 697.400000n V_hig
+ 697.400001n V_hig
+ 697.500000n V_hig
+ 697.500001n V_hig
+ 697.600000n V_hig
+ 697.600001n V_hig
+ 697.700000n V_hig
+ 697.700001n V_hig
+ 697.800000n V_hig
+ 697.800001n V_hig
+ 697.900000n V_hig
+ 697.900001n V_hig
+ 698.000000n V_hig
+ 698.000001n V_hig
+ 698.100000n V_hig
+ 698.100001n V_hig
+ 698.200000n V_hig
+ 698.200001n V_hig
+ 698.300000n V_hig
+ 698.300001n V_hig
+ 698.400000n V_hig
+ 698.400001n V_hig
+ 698.500000n V_hig
+ 698.500001n V_hig
+ 698.600000n V_hig
+ 698.600001n V_hig
+ 698.700000n V_hig
+ 698.700001n V_hig
+ 698.800000n V_hig
+ 698.800001n V_hig
+ 698.900000n V_hig
+ 698.900001n V_hig
+ 699.000000n V_hig
+ 699.000001n V_hig
+ 699.100000n V_hig
+ 699.100001n V_hig
+ 699.200000n V_hig
+ 699.200001n V_hig
+ 699.300000n V_hig
+ 699.300001n V_hig
+ 699.400000n V_hig
+ 699.400001n V_hig
+ 699.500000n V_hig
+ 699.500001n V_hig
+ 699.600000n V_hig
+ 699.600001n V_hig
+ 699.700000n V_hig
+ 699.700001n V_hig
+ 699.800000n V_hig
+ 699.800001n V_hig
+ 699.900000n V_hig
+ 699.900001n V_hig
+ 700.000000n V_hig
+ 700.000001n V_low
+ 700.100000n V_low
+ 700.100001n V_low
+ 700.200000n V_low
+ 700.200001n V_low
+ 700.300000n V_low
+ 700.300001n V_low
+ 700.400000n V_low
+ 700.400001n V_low
+ 700.500000n V_low
+ 700.500001n V_low
+ 700.600000n V_low
+ 700.600001n V_low
+ 700.700000n V_low
+ 700.700001n V_low
+ 700.800000n V_low
+ 700.800001n V_low
+ 700.900000n V_low
+ 700.900001n V_low
+ 701.000000n V_low
+ 701.000001n V_low
+ 701.100000n V_low
+ 701.100001n V_low
+ 701.200000n V_low
+ 701.200001n V_low
+ 701.300000n V_low
+ 701.300001n V_low
+ 701.400000n V_low
+ 701.400001n V_low
+ 701.500000n V_low
+ 701.500001n V_low
+ 701.600000n V_low
+ 701.600001n V_low
+ 701.700000n V_low
+ 701.700001n V_low
+ 701.800000n V_low
+ 701.800001n V_low
+ 701.900000n V_low
+ 701.900001n V_low
+ 702.000000n V_low
+ 702.000001n V_low
+ 702.100000n V_low
+ 702.100001n V_low
+ 702.200000n V_low
+ 702.200001n V_low
+ 702.300000n V_low
+ 702.300001n V_low
+ 702.400000n V_low
+ 702.400001n V_low
+ 702.500000n V_low
+ 702.500001n V_low
+ 702.600000n V_low
+ 702.600001n V_low
+ 702.700000n V_low
+ 702.700001n V_low
+ 702.800000n V_low
+ 702.800001n V_low
+ 702.900000n V_low
+ 702.900001n V_low
+ 703.000000n V_low
+ 703.000001n V_low
+ 703.100000n V_low
+ 703.100001n V_low
+ 703.200000n V_low
+ 703.200001n V_low
+ 703.300000n V_low
+ 703.300001n V_low
+ 703.400000n V_low
+ 703.400001n V_low
+ 703.500000n V_low
+ 703.500001n V_low
+ 703.600000n V_low
+ 703.600001n V_low
+ 703.700000n V_low
+ 703.700001n V_low
+ 703.800000n V_low
+ 703.800001n V_low
+ 703.900000n V_low
+ 703.900001n V_low
+ 704.000000n V_low
+ 704.000001n V_low
+ 704.100000n V_low
+ 704.100001n V_low
+ 704.200000n V_low
+ 704.200001n V_low
+ 704.300000n V_low
+ 704.300001n V_low
+ 704.400000n V_low
+ 704.400001n V_low
+ 704.500000n V_low
+ 704.500001n V_low
+ 704.600000n V_low
+ 704.600001n V_low
+ 704.700000n V_low
+ 704.700001n V_low
+ 704.800000n V_low
+ 704.800001n V_low
+ 704.900000n V_low
+ 704.900001n V_low
+ 705.000000n V_low
+ 705.000001n V_low
+ 705.100000n V_low
+ 705.100001n V_low
+ 705.200000n V_low
+ 705.200001n V_low
+ 705.300000n V_low
+ 705.300001n V_low
+ 705.400000n V_low
+ 705.400001n V_low
+ 705.500000n V_low
+ 705.500001n V_low
+ 705.600000n V_low
+ 705.600001n V_low
+ 705.700000n V_low
+ 705.700001n V_low
+ 705.800000n V_low
+ 705.800001n V_low
+ 705.900000n V_low
+ 705.900001n V_low
+ 706.000000n V_low
+ 706.000001n V_low
+ 706.100000n V_low
+ 706.100001n V_low
+ 706.200000n V_low
+ 706.200001n V_low
+ 706.300000n V_low
+ 706.300001n V_low
+ 706.400000n V_low
+ 706.400001n V_low
+ 706.500000n V_low
+ 706.500001n V_low
+ 706.600000n V_low
+ 706.600001n V_low
+ 706.700000n V_low
+ 706.700001n V_low
+ 706.800000n V_low
+ 706.800001n V_low
+ 706.900000n V_low
+ 706.900001n V_low
+ 707.000000n V_low
+ 707.000001n V_hig
+ 707.100000n V_hig
+ 707.100001n V_hig
+ 707.200000n V_hig
+ 707.200001n V_hig
+ 707.300000n V_hig
+ 707.300001n V_hig
+ 707.400000n V_hig
+ 707.400001n V_hig
+ 707.500000n V_hig
+ 707.500001n V_hig
+ 707.600000n V_hig
+ 707.600001n V_hig
+ 707.700000n V_hig
+ 707.700001n V_hig
+ 707.800000n V_hig
+ 707.800001n V_hig
+ 707.900000n V_hig
+ 707.900001n V_hig
+ 708.000000n V_hig
+ 708.000001n V_low
+ 708.100000n V_low
+ 708.100001n V_low
+ 708.200000n V_low
+ 708.200001n V_low
+ 708.300000n V_low
+ 708.300001n V_low
+ 708.400000n V_low
+ 708.400001n V_low
+ 708.500000n V_low
+ 708.500001n V_low
+ 708.600000n V_low
+ 708.600001n V_low
+ 708.700000n V_low
+ 708.700001n V_low
+ 708.800000n V_low
+ 708.800001n V_low
+ 708.900000n V_low
+ 708.900001n V_low
+ 709.000000n V_low
+ 709.000001n V_low
+ 709.100000n V_low
+ 709.100001n V_low
+ 709.200000n V_low
+ 709.200001n V_low
+ 709.300000n V_low
+ 709.300001n V_low
+ 709.400000n V_low
+ 709.400001n V_low
+ 709.500000n V_low
+ 709.500001n V_low
+ 709.600000n V_low
+ 709.600001n V_low
+ 709.700000n V_low
+ 709.700001n V_low
+ 709.800000n V_low
+ 709.800001n V_low
+ 709.900000n V_low
+ 709.900001n V_low
+ 710.000000n V_low
+ 710.000001n V_hig
+ 710.100000n V_hig
+ 710.100001n V_hig
+ 710.200000n V_hig
+ 710.200001n V_hig
+ 710.300000n V_hig
+ 710.300001n V_hig
+ 710.400000n V_hig
+ 710.400001n V_hig
+ 710.500000n V_hig
+ 710.500001n V_hig
+ 710.600000n V_hig
+ 710.600001n V_hig
+ 710.700000n V_hig
+ 710.700001n V_hig
+ 710.800000n V_hig
+ 710.800001n V_hig
+ 710.900000n V_hig
+ 710.900001n V_hig
+ 711.000000n V_hig
+ 711.000001n V_low
+ 711.100000n V_low
+ 711.100001n V_low
+ 711.200000n V_low
+ 711.200001n V_low
+ 711.300000n V_low
+ 711.300001n V_low
+ 711.400000n V_low
+ 711.400001n V_low
+ 711.500000n V_low
+ 711.500001n V_low
+ 711.600000n V_low
+ 711.600001n V_low
+ 711.700000n V_low
+ 711.700001n V_low
+ 711.800000n V_low
+ 711.800001n V_low
+ 711.900000n V_low
+ 711.900001n V_low
+ 712.000000n V_low
+ 712.000001n V_low
+ 712.100000n V_low
+ 712.100001n V_low
+ 712.200000n V_low
+ 712.200001n V_low
+ 712.300000n V_low
+ 712.300001n V_low
+ 712.400000n V_low
+ 712.400001n V_low
+ 712.500000n V_low
+ 712.500001n V_low
+ 712.600000n V_low
+ 712.600001n V_low
+ 712.700000n V_low
+ 712.700001n V_low
+ 712.800000n V_low
+ 712.800001n V_low
+ 712.900000n V_low
+ 712.900001n V_low
+ 713.000000n V_low
+ 713.000001n V_hig
+ 713.100000n V_hig
+ 713.100001n V_hig
+ 713.200000n V_hig
+ 713.200001n V_hig
+ 713.300000n V_hig
+ 713.300001n V_hig
+ 713.400000n V_hig
+ 713.400001n V_hig
+ 713.500000n V_hig
+ 713.500001n V_hig
+ 713.600000n V_hig
+ 713.600001n V_hig
+ 713.700000n V_hig
+ 713.700001n V_hig
+ 713.800000n V_hig
+ 713.800001n V_hig
+ 713.900000n V_hig
+ 713.900001n V_hig
+ 714.000000n V_hig
+ 714.000001n V_hig
+ 714.100000n V_hig
+ 714.100001n V_hig
+ 714.200000n V_hig
+ 714.200001n V_hig
+ 714.300000n V_hig
+ 714.300001n V_hig
+ 714.400000n V_hig
+ 714.400001n V_hig
+ 714.500000n V_hig
+ 714.500001n V_hig
+ 714.600000n V_hig
+ 714.600001n V_hig
+ 714.700000n V_hig
+ 714.700001n V_hig
+ 714.800000n V_hig
+ 714.800001n V_hig
+ 714.900000n V_hig
+ 714.900001n V_hig
+ 715.000000n V_hig
+ 715.000001n V_hig
+ 715.100000n V_hig
+ 715.100001n V_hig
+ 715.200000n V_hig
+ 715.200001n V_hig
+ 715.300000n V_hig
+ 715.300001n V_hig
+ 715.400000n V_hig
+ 715.400001n V_hig
+ 715.500000n V_hig
+ 715.500001n V_hig
+ 715.600000n V_hig
+ 715.600001n V_hig
+ 715.700000n V_hig
+ 715.700001n V_hig
+ 715.800000n V_hig
+ 715.800001n V_hig
+ 715.900000n V_hig
+ 715.900001n V_hig
+ 716.000000n V_hig
+ 716.000001n V_low
+ 716.100000n V_low
+ 716.100001n V_low
+ 716.200000n V_low
+ 716.200001n V_low
+ 716.300000n V_low
+ 716.300001n V_low
+ 716.400000n V_low
+ 716.400001n V_low
+ 716.500000n V_low
+ 716.500001n V_low
+ 716.600000n V_low
+ 716.600001n V_low
+ 716.700000n V_low
+ 716.700001n V_low
+ 716.800000n V_low
+ 716.800001n V_low
+ 716.900000n V_low
+ 716.900001n V_low
+ 717.000000n V_low
+ 717.000001n V_hig
+ 717.100000n V_hig
+ 717.100001n V_hig
+ 717.200000n V_hig
+ 717.200001n V_hig
+ 717.300000n V_hig
+ 717.300001n V_hig
+ 717.400000n V_hig
+ 717.400001n V_hig
+ 717.500000n V_hig
+ 717.500001n V_hig
+ 717.600000n V_hig
+ 717.600001n V_hig
+ 717.700000n V_hig
+ 717.700001n V_hig
+ 717.800000n V_hig
+ 717.800001n V_hig
+ 717.900000n V_hig
+ 717.900001n V_hig
+ 718.000000n V_hig
+ 718.000001n V_hig
+ 718.100000n V_hig
+ 718.100001n V_hig
+ 718.200000n V_hig
+ 718.200001n V_hig
+ 718.300000n V_hig
+ 718.300001n V_hig
+ 718.400000n V_hig
+ 718.400001n V_hig
+ 718.500000n V_hig
+ 718.500001n V_hig
+ 718.600000n V_hig
+ 718.600001n V_hig
+ 718.700000n V_hig
+ 718.700001n V_hig
+ 718.800000n V_hig
+ 718.800001n V_hig
+ 718.900000n V_hig
+ 718.900001n V_hig
+ 719.000000n V_hig
+ 719.000001n V_hig
+ 719.100000n V_hig
+ 719.100001n V_hig
+ 719.200000n V_hig
+ 719.200001n V_hig
+ 719.300000n V_hig
+ 719.300001n V_hig
+ 719.400000n V_hig
+ 719.400001n V_hig
+ 719.500000n V_hig
+ 719.500001n V_hig
+ 719.600000n V_hig
+ 719.600001n V_hig
+ 719.700000n V_hig
+ 719.700001n V_hig
+ 719.800000n V_hig
+ 719.800001n V_hig
+ 719.900000n V_hig
+ 719.900001n V_hig
+ 720.000000n V_hig
+ 720.000001n V_low
+ 720.100000n V_low
+ 720.100001n V_low
+ 720.200000n V_low
+ 720.200001n V_low
+ 720.300000n V_low
+ 720.300001n V_low
+ 720.400000n V_low
+ 720.400001n V_low
+ 720.500000n V_low
+ 720.500001n V_low
+ 720.600000n V_low
+ 720.600001n V_low
+ 720.700000n V_low
+ 720.700001n V_low
+ 720.800000n V_low
+ 720.800001n V_low
+ 720.900000n V_low
+ 720.900001n V_low
+ 721.000000n V_low
+ 721.000001n V_hig
+ 721.100000n V_hig
+ 721.100001n V_hig
+ 721.200000n V_hig
+ 721.200001n V_hig
+ 721.300000n V_hig
+ 721.300001n V_hig
+ 721.400000n V_hig
+ 721.400001n V_hig
+ 721.500000n V_hig
+ 721.500001n V_hig
+ 721.600000n V_hig
+ 721.600001n V_hig
+ 721.700000n V_hig
+ 721.700001n V_hig
+ 721.800000n V_hig
+ 721.800001n V_hig
+ 721.900000n V_hig
+ 721.900001n V_hig
+ 722.000000n V_hig
+ 722.000001n V_hig
+ 722.100000n V_hig
+ 722.100001n V_hig
+ 722.200000n V_hig
+ 722.200001n V_hig
+ 722.300000n V_hig
+ 722.300001n V_hig
+ 722.400000n V_hig
+ 722.400001n V_hig
+ 722.500000n V_hig
+ 722.500001n V_hig
+ 722.600000n V_hig
+ 722.600001n V_hig
+ 722.700000n V_hig
+ 722.700001n V_hig
+ 722.800000n V_hig
+ 722.800001n V_hig
+ 722.900000n V_hig
+ 722.900001n V_hig
+ 723.000000n V_hig
+ 723.000001n V_low
+ 723.100000n V_low
+ 723.100001n V_low
+ 723.200000n V_low
+ 723.200001n V_low
+ 723.300000n V_low
+ 723.300001n V_low
+ 723.400000n V_low
+ 723.400001n V_low
+ 723.500000n V_low
+ 723.500001n V_low
+ 723.600000n V_low
+ 723.600001n V_low
+ 723.700000n V_low
+ 723.700001n V_low
+ 723.800000n V_low
+ 723.800001n V_low
+ 723.900000n V_low
+ 723.900001n V_low
+ 724.000000n V_low
+ 724.000001n V_hig
+ 724.100000n V_hig
+ 724.100001n V_hig
+ 724.200000n V_hig
+ 724.200001n V_hig
+ 724.300000n V_hig
+ 724.300001n V_hig
+ 724.400000n V_hig
+ 724.400001n V_hig
+ 724.500000n V_hig
+ 724.500001n V_hig
+ 724.600000n V_hig
+ 724.600001n V_hig
+ 724.700000n V_hig
+ 724.700001n V_hig
+ 724.800000n V_hig
+ 724.800001n V_hig
+ 724.900000n V_hig
+ 724.900001n V_hig
+ 725.000000n V_hig
+ 725.000001n V_low
+ 725.100000n V_low
+ 725.100001n V_low
+ 725.200000n V_low
+ 725.200001n V_low
+ 725.300000n V_low
+ 725.300001n V_low
+ 725.400000n V_low
+ 725.400001n V_low
+ 725.500000n V_low
+ 725.500001n V_low
+ 725.600000n V_low
+ 725.600001n V_low
+ 725.700000n V_low
+ 725.700001n V_low
+ 725.800000n V_low
+ 725.800001n V_low
+ 725.900000n V_low
+ 725.900001n V_low
+ 726.000000n V_low
+ 726.000001n V_hig
+ 726.100000n V_hig
+ 726.100001n V_hig
+ 726.200000n V_hig
+ 726.200001n V_hig
+ 726.300000n V_hig
+ 726.300001n V_hig
+ 726.400000n V_hig
+ 726.400001n V_hig
+ 726.500000n V_hig
+ 726.500001n V_hig
+ 726.600000n V_hig
+ 726.600001n V_hig
+ 726.700000n V_hig
+ 726.700001n V_hig
+ 726.800000n V_hig
+ 726.800001n V_hig
+ 726.900000n V_hig
+ 726.900001n V_hig
+ 727.000000n V_hig
+ 727.000001n V_hig
+ 727.100000n V_hig
+ 727.100001n V_hig
+ 727.200000n V_hig
+ 727.200001n V_hig
+ 727.300000n V_hig
+ 727.300001n V_hig
+ 727.400000n V_hig
+ 727.400001n V_hig
+ 727.500000n V_hig
+ 727.500001n V_hig
+ 727.600000n V_hig
+ 727.600001n V_hig
+ 727.700000n V_hig
+ 727.700001n V_hig
+ 727.800000n V_hig
+ 727.800001n V_hig
+ 727.900000n V_hig
+ 727.900001n V_hig
+ 728.000000n V_hig
+ 728.000001n V_hig
+ 728.100000n V_hig
+ 728.100001n V_hig
+ 728.200000n V_hig
+ 728.200001n V_hig
+ 728.300000n V_hig
+ 728.300001n V_hig
+ 728.400000n V_hig
+ 728.400001n V_hig
+ 728.500000n V_hig
+ 728.500001n V_hig
+ 728.600000n V_hig
+ 728.600001n V_hig
+ 728.700000n V_hig
+ 728.700001n V_hig
+ 728.800000n V_hig
+ 728.800001n V_hig
+ 728.900000n V_hig
+ 728.900001n V_hig
+ 729.000000n V_hig
+ 729.000001n V_low
+ 729.100000n V_low
+ 729.100001n V_low
+ 729.200000n V_low
+ 729.200001n V_low
+ 729.300000n V_low
+ 729.300001n V_low
+ 729.400000n V_low
+ 729.400001n V_low
+ 729.500000n V_low
+ 729.500001n V_low
+ 729.600000n V_low
+ 729.600001n V_low
+ 729.700000n V_low
+ 729.700001n V_low
+ 729.800000n V_low
+ 729.800001n V_low
+ 729.900000n V_low
+ 729.900001n V_low
+ 730.000000n V_low
+ 730.000001n V_hig
+ 730.100000n V_hig
+ 730.100001n V_hig
+ 730.200000n V_hig
+ 730.200001n V_hig
+ 730.300000n V_hig
+ 730.300001n V_hig
+ 730.400000n V_hig
+ 730.400001n V_hig
+ 730.500000n V_hig
+ 730.500001n V_hig
+ 730.600000n V_hig
+ 730.600001n V_hig
+ 730.700000n V_hig
+ 730.700001n V_hig
+ 730.800000n V_hig
+ 730.800001n V_hig
+ 730.900000n V_hig
+ 730.900001n V_hig
+ 731.000000n V_hig
+ 731.000001n V_hig
+ 731.100000n V_hig
+ 731.100001n V_hig
+ 731.200000n V_hig
+ 731.200001n V_hig
+ 731.300000n V_hig
+ 731.300001n V_hig
+ 731.400000n V_hig
+ 731.400001n V_hig
+ 731.500000n V_hig
+ 731.500001n V_hig
+ 731.600000n V_hig
+ 731.600001n V_hig
+ 731.700000n V_hig
+ 731.700001n V_hig
+ 731.800000n V_hig
+ 731.800001n V_hig
+ 731.900000n V_hig
+ 731.900001n V_hig
+ 732.000000n V_hig
+ 732.000001n V_hig
+ 732.100000n V_hig
+ 732.100001n V_hig
+ 732.200000n V_hig
+ 732.200001n V_hig
+ 732.300000n V_hig
+ 732.300001n V_hig
+ 732.400000n V_hig
+ 732.400001n V_hig
+ 732.500000n V_hig
+ 732.500001n V_hig
+ 732.600000n V_hig
+ 732.600001n V_hig
+ 732.700000n V_hig
+ 732.700001n V_hig
+ 732.800000n V_hig
+ 732.800001n V_hig
+ 732.900000n V_hig
+ 732.900001n V_hig
+ 733.000000n V_hig
+ 733.000001n V_hig
+ 733.100000n V_hig
+ 733.100001n V_hig
+ 733.200000n V_hig
+ 733.200001n V_hig
+ 733.300000n V_hig
+ 733.300001n V_hig
+ 733.400000n V_hig
+ 733.400001n V_hig
+ 733.500000n V_hig
+ 733.500001n V_hig
+ 733.600000n V_hig
+ 733.600001n V_hig
+ 733.700000n V_hig
+ 733.700001n V_hig
+ 733.800000n V_hig
+ 733.800001n V_hig
+ 733.900000n V_hig
+ 733.900001n V_hig
+ 734.000000n V_hig
+ 734.000001n V_hig
+ 734.100000n V_hig
+ 734.100001n V_hig
+ 734.200000n V_hig
+ 734.200001n V_hig
+ 734.300000n V_hig
+ 734.300001n V_hig
+ 734.400000n V_hig
+ 734.400001n V_hig
+ 734.500000n V_hig
+ 734.500001n V_hig
+ 734.600000n V_hig
+ 734.600001n V_hig
+ 734.700000n V_hig
+ 734.700001n V_hig
+ 734.800000n V_hig
+ 734.800001n V_hig
+ 734.900000n V_hig
+ 734.900001n V_hig
+ 735.000000n V_hig
+ 735.000001n V_hig
+ 735.100000n V_hig
+ 735.100001n V_hig
+ 735.200000n V_hig
+ 735.200001n V_hig
+ 735.300000n V_hig
+ 735.300001n V_hig
+ 735.400000n V_hig
+ 735.400001n V_hig
+ 735.500000n V_hig
+ 735.500001n V_hig
+ 735.600000n V_hig
+ 735.600001n V_hig
+ 735.700000n V_hig
+ 735.700001n V_hig
+ 735.800000n V_hig
+ 735.800001n V_hig
+ 735.900000n V_hig
+ 735.900001n V_hig
+ 736.000000n V_hig
+ 736.000001n V_hig
+ 736.100000n V_hig
+ 736.100001n V_hig
+ 736.200000n V_hig
+ 736.200001n V_hig
+ 736.300000n V_hig
+ 736.300001n V_hig
+ 736.400000n V_hig
+ 736.400001n V_hig
+ 736.500000n V_hig
+ 736.500001n V_hig
+ 736.600000n V_hig
+ 736.600001n V_hig
+ 736.700000n V_hig
+ 736.700001n V_hig
+ 736.800000n V_hig
+ 736.800001n V_hig
+ 736.900000n V_hig
+ 736.900001n V_hig
+ 737.000000n V_hig
+ 737.000001n V_hig
+ 737.100000n V_hig
+ 737.100001n V_hig
+ 737.200000n V_hig
+ 737.200001n V_hig
+ 737.300000n V_hig
+ 737.300001n V_hig
+ 737.400000n V_hig
+ 737.400001n V_hig
+ 737.500000n V_hig
+ 737.500001n V_hig
+ 737.600000n V_hig
+ 737.600001n V_hig
+ 737.700000n V_hig
+ 737.700001n V_hig
+ 737.800000n V_hig
+ 737.800001n V_hig
+ 737.900000n V_hig
+ 737.900001n V_hig
+ 738.000000n V_hig
+ 738.000001n V_hig
+ 738.100000n V_hig
+ 738.100001n V_hig
+ 738.200000n V_hig
+ 738.200001n V_hig
+ 738.300000n V_hig
+ 738.300001n V_hig
+ 738.400000n V_hig
+ 738.400001n V_hig
+ 738.500000n V_hig
+ 738.500001n V_hig
+ 738.600000n V_hig
+ 738.600001n V_hig
+ 738.700000n V_hig
+ 738.700001n V_hig
+ 738.800000n V_hig
+ 738.800001n V_hig
+ 738.900000n V_hig
+ 738.900001n V_hig
+ 739.000000n V_hig
+ 739.000001n V_hig
+ 739.100000n V_hig
+ 739.100001n V_hig
+ 739.200000n V_hig
+ 739.200001n V_hig
+ 739.300000n V_hig
+ 739.300001n V_hig
+ 739.400000n V_hig
+ 739.400001n V_hig
+ 739.500000n V_hig
+ 739.500001n V_hig
+ 739.600000n V_hig
+ 739.600001n V_hig
+ 739.700000n V_hig
+ 739.700001n V_hig
+ 739.800000n V_hig
+ 739.800001n V_hig
+ 739.900000n V_hig
+ 739.900001n V_hig
+ 740.000000n V_hig
+ 740.000001n V_hig
+ 740.100000n V_hig
+ 740.100001n V_hig
+ 740.200000n V_hig
+ 740.200001n V_hig
+ 740.300000n V_hig
+ 740.300001n V_hig
+ 740.400000n V_hig
+ 740.400001n V_hig
+ 740.500000n V_hig
+ 740.500001n V_hig
+ 740.600000n V_hig
+ 740.600001n V_hig
+ 740.700000n V_hig
+ 740.700001n V_hig
+ 740.800000n V_hig
+ 740.800001n V_hig
+ 740.900000n V_hig
+ 740.900001n V_hig
+ 741.000000n V_hig
+ 741.000001n V_hig
+ 741.100000n V_hig
+ 741.100001n V_hig
+ 741.200000n V_hig
+ 741.200001n V_hig
+ 741.300000n V_hig
+ 741.300001n V_hig
+ 741.400000n V_hig
+ 741.400001n V_hig
+ 741.500000n V_hig
+ 741.500001n V_hig
+ 741.600000n V_hig
+ 741.600001n V_hig
+ 741.700000n V_hig
+ 741.700001n V_hig
+ 741.800000n V_hig
+ 741.800001n V_hig
+ 741.900000n V_hig
+ 741.900001n V_hig
+ 742.000000n V_hig
+ 742.000001n V_low
+ 742.100000n V_low
+ 742.100001n V_low
+ 742.200000n V_low
+ 742.200001n V_low
+ 742.300000n V_low
+ 742.300001n V_low
+ 742.400000n V_low
+ 742.400001n V_low
+ 742.500000n V_low
+ 742.500001n V_low
+ 742.600000n V_low
+ 742.600001n V_low
+ 742.700000n V_low
+ 742.700001n V_low
+ 742.800000n V_low
+ 742.800001n V_low
+ 742.900000n V_low
+ 742.900001n V_low
+ 743.000000n V_low
+ 743.000001n V_hig
+ 743.100000n V_hig
+ 743.100001n V_hig
+ 743.200000n V_hig
+ 743.200001n V_hig
+ 743.300000n V_hig
+ 743.300001n V_hig
+ 743.400000n V_hig
+ 743.400001n V_hig
+ 743.500000n V_hig
+ 743.500001n V_hig
+ 743.600000n V_hig
+ 743.600001n V_hig
+ 743.700000n V_hig
+ 743.700001n V_hig
+ 743.800000n V_hig
+ 743.800001n V_hig
+ 743.900000n V_hig
+ 743.900001n V_hig
+ 744.000000n V_hig
+ 744.000001n V_hig
+ 744.100000n V_hig
+ 744.100001n V_hig
+ 744.200000n V_hig
+ 744.200001n V_hig
+ 744.300000n V_hig
+ 744.300001n V_hig
+ 744.400000n V_hig
+ 744.400001n V_hig
+ 744.500000n V_hig
+ 744.500001n V_hig
+ 744.600000n V_hig
+ 744.600001n V_hig
+ 744.700000n V_hig
+ 744.700001n V_hig
+ 744.800000n V_hig
+ 744.800001n V_hig
+ 744.900000n V_hig
+ 744.900001n V_hig
+ 745.000000n V_hig
+ 745.000001n V_low
+ 745.100000n V_low
+ 745.100001n V_low
+ 745.200000n V_low
+ 745.200001n V_low
+ 745.300000n V_low
+ 745.300001n V_low
+ 745.400000n V_low
+ 745.400001n V_low
+ 745.500000n V_low
+ 745.500001n V_low
+ 745.600000n V_low
+ 745.600001n V_low
+ 745.700000n V_low
+ 745.700001n V_low
+ 745.800000n V_low
+ 745.800001n V_low
+ 745.900000n V_low
+ 745.900001n V_low
+ 746.000000n V_low
+ 746.000001n V_low
+ 746.100000n V_low
+ 746.100001n V_low
+ 746.200000n V_low
+ 746.200001n V_low
+ 746.300000n V_low
+ 746.300001n V_low
+ 746.400000n V_low
+ 746.400001n V_low
+ 746.500000n V_low
+ 746.500001n V_low
+ 746.600000n V_low
+ 746.600001n V_low
+ 746.700000n V_low
+ 746.700001n V_low
+ 746.800000n V_low
+ 746.800001n V_low
+ 746.900000n V_low
+ 746.900001n V_low
+ 747.000000n V_low
+ 747.000001n V_low
+ 747.100000n V_low
+ 747.100001n V_low
+ 747.200000n V_low
+ 747.200001n V_low
+ 747.300000n V_low
+ 747.300001n V_low
+ 747.400000n V_low
+ 747.400001n V_low
+ 747.500000n V_low
+ 747.500001n V_low
+ 747.600000n V_low
+ 747.600001n V_low
+ 747.700000n V_low
+ 747.700001n V_low
+ 747.800000n V_low
+ 747.800001n V_low
+ 747.900000n V_low
+ 747.900001n V_low
+ 748.000000n V_low
+ 748.000001n V_low
+ 748.100000n V_low
+ 748.100001n V_low
+ 748.200000n V_low
+ 748.200001n V_low
+ 748.300000n V_low
+ 748.300001n V_low
+ 748.400000n V_low
+ 748.400001n V_low
+ 748.500000n V_low
+ 748.500001n V_low
+ 748.600000n V_low
+ 748.600001n V_low
+ 748.700000n V_low
+ 748.700001n V_low
+ 748.800000n V_low
+ 748.800001n V_low
+ 748.900000n V_low
+ 748.900001n V_low
+ 749.000000n V_low
+ 749.000001n V_low
+ 749.100000n V_low
+ 749.100001n V_low
+ 749.200000n V_low
+ 749.200001n V_low
+ 749.300000n V_low
+ 749.300001n V_low
+ 749.400000n V_low
+ 749.400001n V_low
+ 749.500000n V_low
+ 749.500001n V_low
+ 749.600000n V_low
+ 749.600001n V_low
+ 749.700000n V_low
+ 749.700001n V_low
+ 749.800000n V_low
+ 749.800001n V_low
+ 749.900000n V_low
+ 749.900001n V_low
+ 750.000000n V_low
+ 750.000001n V_hig
+ 750.100000n V_hig
+ 750.100001n V_hig
+ 750.200000n V_hig
+ 750.200001n V_hig
+ 750.300000n V_hig
+ 750.300001n V_hig
+ 750.400000n V_hig
+ 750.400001n V_hig
+ 750.500000n V_hig
+ 750.500001n V_hig
+ 750.600000n V_hig
+ 750.600001n V_hig
+ 750.700000n V_hig
+ 750.700001n V_hig
+ 750.800000n V_hig
+ 750.800001n V_hig
+ 750.900000n V_hig
+ 750.900001n V_hig
+ 751.000000n V_hig
+ 751.000001n V_hig
+ 751.100000n V_hig
+ 751.100001n V_hig
+ 751.200000n V_hig
+ 751.200001n V_hig
+ 751.300000n V_hig
+ 751.300001n V_hig
+ 751.400000n V_hig
+ 751.400001n V_hig
+ 751.500000n V_hig
+ 751.500001n V_hig
+ 751.600000n V_hig
+ 751.600001n V_hig
+ 751.700000n V_hig
+ 751.700001n V_hig
+ 751.800000n V_hig
+ 751.800001n V_hig
+ 751.900000n V_hig
+ 751.900001n V_hig
+ 752.000000n V_hig
+ 752.000001n V_low
+ 752.100000n V_low
+ 752.100001n V_low
+ 752.200000n V_low
+ 752.200001n V_low
+ 752.300000n V_low
+ 752.300001n V_low
+ 752.400000n V_low
+ 752.400001n V_low
+ 752.500000n V_low
+ 752.500001n V_low
+ 752.600000n V_low
+ 752.600001n V_low
+ 752.700000n V_low
+ 752.700001n V_low
+ 752.800000n V_low
+ 752.800001n V_low
+ 752.900000n V_low
+ 752.900001n V_low
+ 753.000000n V_low
+ 753.000001n V_low
+ 753.100000n V_low
+ 753.100001n V_low
+ 753.200000n V_low
+ 753.200001n V_low
+ 753.300000n V_low
+ 753.300001n V_low
+ 753.400000n V_low
+ 753.400001n V_low
+ 753.500000n V_low
+ 753.500001n V_low
+ 753.600000n V_low
+ 753.600001n V_low
+ 753.700000n V_low
+ 753.700001n V_low
+ 753.800000n V_low
+ 753.800001n V_low
+ 753.900000n V_low
+ 753.900001n V_low
+ 754.000000n V_low
+ 754.000001n V_hig
+ 754.100000n V_hig
+ 754.100001n V_hig
+ 754.200000n V_hig
+ 754.200001n V_hig
+ 754.300000n V_hig
+ 754.300001n V_hig
+ 754.400000n V_hig
+ 754.400001n V_hig
+ 754.500000n V_hig
+ 754.500001n V_hig
+ 754.600000n V_hig
+ 754.600001n V_hig
+ 754.700000n V_hig
+ 754.700001n V_hig
+ 754.800000n V_hig
+ 754.800001n V_hig
+ 754.900000n V_hig
+ 754.900001n V_hig
+ 755.000000n V_hig
+ 755.000001n V_low
+ 755.100000n V_low
+ 755.100001n V_low
+ 755.200000n V_low
+ 755.200001n V_low
+ 755.300000n V_low
+ 755.300001n V_low
+ 755.400000n V_low
+ 755.400001n V_low
+ 755.500000n V_low
+ 755.500001n V_low
+ 755.600000n V_low
+ 755.600001n V_low
+ 755.700000n V_low
+ 755.700001n V_low
+ 755.800000n V_low
+ 755.800001n V_low
+ 755.900000n V_low
+ 755.900001n V_low
+ 756.000000n V_low
+ 756.000001n V_hig
+ 756.100000n V_hig
+ 756.100001n V_hig
+ 756.200000n V_hig
+ 756.200001n V_hig
+ 756.300000n V_hig
+ 756.300001n V_hig
+ 756.400000n V_hig
+ 756.400001n V_hig
+ 756.500000n V_hig
+ 756.500001n V_hig
+ 756.600000n V_hig
+ 756.600001n V_hig
+ 756.700000n V_hig
+ 756.700001n V_hig
+ 756.800000n V_hig
+ 756.800001n V_hig
+ 756.900000n V_hig
+ 756.900001n V_hig
+ 757.000000n V_hig
+ 757.000001n V_low
+ 757.100000n V_low
+ 757.100001n V_low
+ 757.200000n V_low
+ 757.200001n V_low
+ 757.300000n V_low
+ 757.300001n V_low
+ 757.400000n V_low
+ 757.400001n V_low
+ 757.500000n V_low
+ 757.500001n V_low
+ 757.600000n V_low
+ 757.600001n V_low
+ 757.700000n V_low
+ 757.700001n V_low
+ 757.800000n V_low
+ 757.800001n V_low
+ 757.900000n V_low
+ 757.900001n V_low
+ 758.000000n V_low
+ 758.000001n V_hig
+ 758.100000n V_hig
+ 758.100001n V_hig
+ 758.200000n V_hig
+ 758.200001n V_hig
+ 758.300000n V_hig
+ 758.300001n V_hig
+ 758.400000n V_hig
+ 758.400001n V_hig
+ 758.500000n V_hig
+ 758.500001n V_hig
+ 758.600000n V_hig
+ 758.600001n V_hig
+ 758.700000n V_hig
+ 758.700001n V_hig
+ 758.800000n V_hig
+ 758.800001n V_hig
+ 758.900000n V_hig
+ 758.900001n V_hig
+ 759.000000n V_hig
+ 759.000001n V_low
+ 759.100000n V_low
+ 759.100001n V_low
+ 759.200000n V_low
+ 759.200001n V_low
+ 759.300000n V_low
+ 759.300001n V_low
+ 759.400000n V_low
+ 759.400001n V_low
+ 759.500000n V_low
+ 759.500001n V_low
+ 759.600000n V_low
+ 759.600001n V_low
+ 759.700000n V_low
+ 759.700001n V_low
+ 759.800000n V_low
+ 759.800001n V_low
+ 759.900000n V_low
+ 759.900001n V_low
+ 760.000000n V_low
+ 760.000001n V_low
+ 760.100000n V_low
+ 760.100001n V_low
+ 760.200000n V_low
+ 760.200001n V_low
+ 760.300000n V_low
+ 760.300001n V_low
+ 760.400000n V_low
+ 760.400001n V_low
+ 760.500000n V_low
+ 760.500001n V_low
+ 760.600000n V_low
+ 760.600001n V_low
+ 760.700000n V_low
+ 760.700001n V_low
+ 760.800000n V_low
+ 760.800001n V_low
+ 760.900000n V_low
+ 760.900001n V_low
+ 761.000000n V_low
+ 761.000001n V_low
+ 761.100000n V_low
+ 761.100001n V_low
+ 761.200000n V_low
+ 761.200001n V_low
+ 761.300000n V_low
+ 761.300001n V_low
+ 761.400000n V_low
+ 761.400001n V_low
+ 761.500000n V_low
+ 761.500001n V_low
+ 761.600000n V_low
+ 761.600001n V_low
+ 761.700000n V_low
+ 761.700001n V_low
+ 761.800000n V_low
+ 761.800001n V_low
+ 761.900000n V_low
+ 761.900001n V_low
+ 762.000000n V_low
+ 762.000001n V_low
+ 762.100000n V_low
+ 762.100001n V_low
+ 762.200000n V_low
+ 762.200001n V_low
+ 762.300000n V_low
+ 762.300001n V_low
+ 762.400000n V_low
+ 762.400001n V_low
+ 762.500000n V_low
+ 762.500001n V_low
+ 762.600000n V_low
+ 762.600001n V_low
+ 762.700000n V_low
+ 762.700001n V_low
+ 762.800000n V_low
+ 762.800001n V_low
+ 762.900000n V_low
+ 762.900001n V_low
+ 763.000000n V_low
+ 763.000001n V_low
+ 763.100000n V_low
+ 763.100001n V_low
+ 763.200000n V_low
+ 763.200001n V_low
+ 763.300000n V_low
+ 763.300001n V_low
+ 763.400000n V_low
+ 763.400001n V_low
+ 763.500000n V_low
+ 763.500001n V_low
+ 763.600000n V_low
+ 763.600001n V_low
+ 763.700000n V_low
+ 763.700001n V_low
+ 763.800000n V_low
+ 763.800001n V_low
+ 763.900000n V_low
+ 763.900001n V_low
+ 764.000000n V_low
+ 764.000001n V_hig
+ 764.100000n V_hig
+ 764.100001n V_hig
+ 764.200000n V_hig
+ 764.200001n V_hig
+ 764.300000n V_hig
+ 764.300001n V_hig
+ 764.400000n V_hig
+ 764.400001n V_hig
+ 764.500000n V_hig
+ 764.500001n V_hig
+ 764.600000n V_hig
+ 764.600001n V_hig
+ 764.700000n V_hig
+ 764.700001n V_hig
+ 764.800000n V_hig
+ 764.800001n V_hig
+ 764.900000n V_hig
+ 764.900001n V_hig
+ 765.000000n V_hig
+ 765.000001n V_hig
+ 765.100000n V_hig
+ 765.100001n V_hig
+ 765.200000n V_hig
+ 765.200001n V_hig
+ 765.300000n V_hig
+ 765.300001n V_hig
+ 765.400000n V_hig
+ 765.400001n V_hig
+ 765.500000n V_hig
+ 765.500001n V_hig
+ 765.600000n V_hig
+ 765.600001n V_hig
+ 765.700000n V_hig
+ 765.700001n V_hig
+ 765.800000n V_hig
+ 765.800001n V_hig
+ 765.900000n V_hig
+ 765.900001n V_hig
+ 766.000000n V_hig
+ 766.000001n V_hig
+ 766.100000n V_hig
+ 766.100001n V_hig
+ 766.200000n V_hig
+ 766.200001n V_hig
+ 766.300000n V_hig
+ 766.300001n V_hig
+ 766.400000n V_hig
+ 766.400001n V_hig
+ 766.500000n V_hig
+ 766.500001n V_hig
+ 766.600000n V_hig
+ 766.600001n V_hig
+ 766.700000n V_hig
+ 766.700001n V_hig
+ 766.800000n V_hig
+ 766.800001n V_hig
+ 766.900000n V_hig
+ 766.900001n V_hig
+ 767.000000n V_hig
+ 767.000001n V_low
+ 767.100000n V_low
+ 767.100001n V_low
+ 767.200000n V_low
+ 767.200001n V_low
+ 767.300000n V_low
+ 767.300001n V_low
+ 767.400000n V_low
+ 767.400001n V_low
+ 767.500000n V_low
+ 767.500001n V_low
+ 767.600000n V_low
+ 767.600001n V_low
+ 767.700000n V_low
+ 767.700001n V_low
+ 767.800000n V_low
+ 767.800001n V_low
+ 767.900000n V_low
+ 767.900001n V_low
+ 768.000000n V_low
+ 768.000001n V_hig
+ 768.100000n V_hig
+ 768.100001n V_hig
+ 768.200000n V_hig
+ 768.200001n V_hig
+ 768.300000n V_hig
+ 768.300001n V_hig
+ 768.400000n V_hig
+ 768.400001n V_hig
+ 768.500000n V_hig
+ 768.500001n V_hig
+ 768.600000n V_hig
+ 768.600001n V_hig
+ 768.700000n V_hig
+ 768.700001n V_hig
+ 768.800000n V_hig
+ 768.800001n V_hig
+ 768.900000n V_hig
+ 768.900001n V_hig
+ 769.000000n V_hig
+ 769.000001n V_hig
+ 769.100000n V_hig
+ 769.100001n V_hig
+ 769.200000n V_hig
+ 769.200001n V_hig
+ 769.300000n V_hig
+ 769.300001n V_hig
+ 769.400000n V_hig
+ 769.400001n V_hig
+ 769.500000n V_hig
+ 769.500001n V_hig
+ 769.600000n V_hig
+ 769.600001n V_hig
+ 769.700000n V_hig
+ 769.700001n V_hig
+ 769.800000n V_hig
+ 769.800001n V_hig
+ 769.900000n V_hig
+ 769.900001n V_hig
+ 770.000000n V_hig
+ 770.000001n V_hig
+ 770.100000n V_hig
+ 770.100001n V_hig
+ 770.200000n V_hig
+ 770.200001n V_hig
+ 770.300000n V_hig
+ 770.300001n V_hig
+ 770.400000n V_hig
+ 770.400001n V_hig
+ 770.500000n V_hig
+ 770.500001n V_hig
+ 770.600000n V_hig
+ 770.600001n V_hig
+ 770.700000n V_hig
+ 770.700001n V_hig
+ 770.800000n V_hig
+ 770.800001n V_hig
+ 770.900000n V_hig
+ 770.900001n V_hig
+ 771.000000n V_hig
+ 771.000001n V_hig
+ 771.100000n V_hig
+ 771.100001n V_hig
+ 771.200000n V_hig
+ 771.200001n V_hig
+ 771.300000n V_hig
+ 771.300001n V_hig
+ 771.400000n V_hig
+ 771.400001n V_hig
+ 771.500000n V_hig
+ 771.500001n V_hig
+ 771.600000n V_hig
+ 771.600001n V_hig
+ 771.700000n V_hig
+ 771.700001n V_hig
+ 771.800000n V_hig
+ 771.800001n V_hig
+ 771.900000n V_hig
+ 771.900001n V_hig
+ 772.000000n V_hig
+ 772.000001n V_hig
+ 772.100000n V_hig
+ 772.100001n V_hig
+ 772.200000n V_hig
+ 772.200001n V_hig
+ 772.300000n V_hig
+ 772.300001n V_hig
+ 772.400000n V_hig
+ 772.400001n V_hig
+ 772.500000n V_hig
+ 772.500001n V_hig
+ 772.600000n V_hig
+ 772.600001n V_hig
+ 772.700000n V_hig
+ 772.700001n V_hig
+ 772.800000n V_hig
+ 772.800001n V_hig
+ 772.900000n V_hig
+ 772.900001n V_hig
+ 773.000000n V_hig
+ 773.000001n V_low
+ 773.100000n V_low
+ 773.100001n V_low
+ 773.200000n V_low
+ 773.200001n V_low
+ 773.300000n V_low
+ 773.300001n V_low
+ 773.400000n V_low
+ 773.400001n V_low
+ 773.500000n V_low
+ 773.500001n V_low
+ 773.600000n V_low
+ 773.600001n V_low
+ 773.700000n V_low
+ 773.700001n V_low
+ 773.800000n V_low
+ 773.800001n V_low
+ 773.900000n V_low
+ 773.900001n V_low
+ 774.000000n V_low
+ 774.000001n V_low
+ 774.100000n V_low
+ 774.100001n V_low
+ 774.200000n V_low
+ 774.200001n V_low
+ 774.300000n V_low
+ 774.300001n V_low
+ 774.400000n V_low
+ 774.400001n V_low
+ 774.500000n V_low
+ 774.500001n V_low
+ 774.600000n V_low
+ 774.600001n V_low
+ 774.700000n V_low
+ 774.700001n V_low
+ 774.800000n V_low
+ 774.800001n V_low
+ 774.900000n V_low
+ 774.900001n V_low
+ 775.000000n V_low
+ 775.000001n V_hig
+ 775.100000n V_hig
+ 775.100001n V_hig
+ 775.200000n V_hig
+ 775.200001n V_hig
+ 775.300000n V_hig
+ 775.300001n V_hig
+ 775.400000n V_hig
+ 775.400001n V_hig
+ 775.500000n V_hig
+ 775.500001n V_hig
+ 775.600000n V_hig
+ 775.600001n V_hig
+ 775.700000n V_hig
+ 775.700001n V_hig
+ 775.800000n V_hig
+ 775.800001n V_hig
+ 775.900000n V_hig
+ 775.900001n V_hig
+ 776.000000n V_hig
+ 776.000001n V_low
+ 776.100000n V_low
+ 776.100001n V_low
+ 776.200000n V_low
+ 776.200001n V_low
+ 776.300000n V_low
+ 776.300001n V_low
+ 776.400000n V_low
+ 776.400001n V_low
+ 776.500000n V_low
+ 776.500001n V_low
+ 776.600000n V_low
+ 776.600001n V_low
+ 776.700000n V_low
+ 776.700001n V_low
+ 776.800000n V_low
+ 776.800001n V_low
+ 776.900000n V_low
+ 776.900001n V_low
+ 777.000000n V_low
+ 777.000001n V_low
+ 777.100000n V_low
+ 777.100001n V_low
+ 777.200000n V_low
+ 777.200001n V_low
+ 777.300000n V_low
+ 777.300001n V_low
+ 777.400000n V_low
+ 777.400001n V_low
+ 777.500000n V_low
+ 777.500001n V_low
+ 777.600000n V_low
+ 777.600001n V_low
+ 777.700000n V_low
+ 777.700001n V_low
+ 777.800000n V_low
+ 777.800001n V_low
+ 777.900000n V_low
+ 777.900001n V_low
+ 778.000000n V_low
+ 778.000001n V_hig
+ 778.100000n V_hig
+ 778.100001n V_hig
+ 778.200000n V_hig
+ 778.200001n V_hig
+ 778.300000n V_hig
+ 778.300001n V_hig
+ 778.400000n V_hig
+ 778.400001n V_hig
+ 778.500000n V_hig
+ 778.500001n V_hig
+ 778.600000n V_hig
+ 778.600001n V_hig
+ 778.700000n V_hig
+ 778.700001n V_hig
+ 778.800000n V_hig
+ 778.800001n V_hig
+ 778.900000n V_hig
+ 778.900001n V_hig
+ 779.000000n V_hig
+ 779.000001n V_hig
+ 779.100000n V_hig
+ 779.100001n V_hig
+ 779.200000n V_hig
+ 779.200001n V_hig
+ 779.300000n V_hig
+ 779.300001n V_hig
+ 779.400000n V_hig
+ 779.400001n V_hig
+ 779.500000n V_hig
+ 779.500001n V_hig
+ 779.600000n V_hig
+ 779.600001n V_hig
+ 779.700000n V_hig
+ 779.700001n V_hig
+ 779.800000n V_hig
+ 779.800001n V_hig
+ 779.900000n V_hig
+ 779.900001n V_hig
+ 780.000000n V_hig
+ 780.000001n V_hig
+ 780.100000n V_hig
+ 780.100001n V_hig
+ 780.200000n V_hig
+ 780.200001n V_hig
+ 780.300000n V_hig
+ 780.300001n V_hig
+ 780.400000n V_hig
+ 780.400001n V_hig
+ 780.500000n V_hig
+ 780.500001n V_hig
+ 780.600000n V_hig
+ 780.600001n V_hig
+ 780.700000n V_hig
+ 780.700001n V_hig
+ 780.800000n V_hig
+ 780.800001n V_hig
+ 780.900000n V_hig
+ 780.900001n V_hig
+ 781.000000n V_hig
+ 781.000001n V_hig
+ 781.100000n V_hig
+ 781.100001n V_hig
+ 781.200000n V_hig
+ 781.200001n V_hig
+ 781.300000n V_hig
+ 781.300001n V_hig
+ 781.400000n V_hig
+ 781.400001n V_hig
+ 781.500000n V_hig
+ 781.500001n V_hig
+ 781.600000n V_hig
+ 781.600001n V_hig
+ 781.700000n V_hig
+ 781.700001n V_hig
+ 781.800000n V_hig
+ 781.800001n V_hig
+ 781.900000n V_hig
+ 781.900001n V_hig
+ 782.000000n V_hig
+ 782.000001n V_low
+ 782.100000n V_low
+ 782.100001n V_low
+ 782.200000n V_low
+ 782.200001n V_low
+ 782.300000n V_low
+ 782.300001n V_low
+ 782.400000n V_low
+ 782.400001n V_low
+ 782.500000n V_low
+ 782.500001n V_low
+ 782.600000n V_low
+ 782.600001n V_low
+ 782.700000n V_low
+ 782.700001n V_low
+ 782.800000n V_low
+ 782.800001n V_low
+ 782.900000n V_low
+ 782.900001n V_low
+ 783.000000n V_low
+ 783.000001n V_hig
+ 783.100000n V_hig
+ 783.100001n V_hig
+ 783.200000n V_hig
+ 783.200001n V_hig
+ 783.300000n V_hig
+ 783.300001n V_hig
+ 783.400000n V_hig
+ 783.400001n V_hig
+ 783.500000n V_hig
+ 783.500001n V_hig
+ 783.600000n V_hig
+ 783.600001n V_hig
+ 783.700000n V_hig
+ 783.700001n V_hig
+ 783.800000n V_hig
+ 783.800001n V_hig
+ 783.900000n V_hig
+ 783.900001n V_hig
+ 784.000000n V_hig
+ 784.000001n V_hig
+ 784.100000n V_hig
+ 784.100001n V_hig
+ 784.200000n V_hig
+ 784.200001n V_hig
+ 784.300000n V_hig
+ 784.300001n V_hig
+ 784.400000n V_hig
+ 784.400001n V_hig
+ 784.500000n V_hig
+ 784.500001n V_hig
+ 784.600000n V_hig
+ 784.600001n V_hig
+ 784.700000n V_hig
+ 784.700001n V_hig
+ 784.800000n V_hig
+ 784.800001n V_hig
+ 784.900000n V_hig
+ 784.900001n V_hig
+ 785.000000n V_hig
+ 785.000001n V_hig
+ 785.100000n V_hig
+ 785.100001n V_hig
+ 785.200000n V_hig
+ 785.200001n V_hig
+ 785.300000n V_hig
+ 785.300001n V_hig
+ 785.400000n V_hig
+ 785.400001n V_hig
+ 785.500000n V_hig
+ 785.500001n V_hig
+ 785.600000n V_hig
+ 785.600001n V_hig
+ 785.700000n V_hig
+ 785.700001n V_hig
+ 785.800000n V_hig
+ 785.800001n V_hig
+ 785.900000n V_hig
+ 785.900001n V_hig
+ 786.000000n V_hig
+ 786.000001n V_hig
+ 786.100000n V_hig
+ 786.100001n V_hig
+ 786.200000n V_hig
+ 786.200001n V_hig
+ 786.300000n V_hig
+ 786.300001n V_hig
+ 786.400000n V_hig
+ 786.400001n V_hig
+ 786.500000n V_hig
+ 786.500001n V_hig
+ 786.600000n V_hig
+ 786.600001n V_hig
+ 786.700000n V_hig
+ 786.700001n V_hig
+ 786.800000n V_hig
+ 786.800001n V_hig
+ 786.900000n V_hig
+ 786.900001n V_hig
+ 787.000000n V_hig
+ 787.000001n V_hig
+ 787.100000n V_hig
+ 787.100001n V_hig
+ 787.200000n V_hig
+ 787.200001n V_hig
+ 787.300000n V_hig
+ 787.300001n V_hig
+ 787.400000n V_hig
+ 787.400001n V_hig
+ 787.500000n V_hig
+ 787.500001n V_hig
+ 787.600000n V_hig
+ 787.600001n V_hig
+ 787.700000n V_hig
+ 787.700001n V_hig
+ 787.800000n V_hig
+ 787.800001n V_hig
+ 787.900000n V_hig
+ 787.900001n V_hig
+ 788.000000n V_hig
+ 788.000001n V_hig
+ 788.100000n V_hig
+ 788.100001n V_hig
+ 788.200000n V_hig
+ 788.200001n V_hig
+ 788.300000n V_hig
+ 788.300001n V_hig
+ 788.400000n V_hig
+ 788.400001n V_hig
+ 788.500000n V_hig
+ 788.500001n V_hig
+ 788.600000n V_hig
+ 788.600001n V_hig
+ 788.700000n V_hig
+ 788.700001n V_hig
+ 788.800000n V_hig
+ 788.800001n V_hig
+ 788.900000n V_hig
+ 788.900001n V_hig
+ 789.000000n V_hig
+ 789.000001n V_low
+ 789.100000n V_low
+ 789.100001n V_low
+ 789.200000n V_low
+ 789.200001n V_low
+ 789.300000n V_low
+ 789.300001n V_low
+ 789.400000n V_low
+ 789.400001n V_low
+ 789.500000n V_low
+ 789.500001n V_low
+ 789.600000n V_low
+ 789.600001n V_low
+ 789.700000n V_low
+ 789.700001n V_low
+ 789.800000n V_low
+ 789.800001n V_low
+ 789.900000n V_low
+ 789.900001n V_low
+ 790.000000n V_low
+ 790.000001n V_low
+ 790.100000n V_low
+ 790.100001n V_low
+ 790.200000n V_low
+ 790.200001n V_low
+ 790.300000n V_low
+ 790.300001n V_low
+ 790.400000n V_low
+ 790.400001n V_low
+ 790.500000n V_low
+ 790.500001n V_low
+ 790.600000n V_low
+ 790.600001n V_low
+ 790.700000n V_low
+ 790.700001n V_low
+ 790.800000n V_low
+ 790.800001n V_low
+ 790.900000n V_low
+ 790.900001n V_low
+ 791.000000n V_low
+ 791.000001n V_low
+ 791.100000n V_low
+ 791.100001n V_low
+ 791.200000n V_low
+ 791.200001n V_low
+ 791.300000n V_low
+ 791.300001n V_low
+ 791.400000n V_low
+ 791.400001n V_low
+ 791.500000n V_low
+ 791.500001n V_low
+ 791.600000n V_low
+ 791.600001n V_low
+ 791.700000n V_low
+ 791.700001n V_low
+ 791.800000n V_low
+ 791.800001n V_low
+ 791.900000n V_low
+ 791.900001n V_low
+ 792.000000n V_low
+ 792.000001n V_low
+ 792.100000n V_low
+ 792.100001n V_low
+ 792.200000n V_low
+ 792.200001n V_low
+ 792.300000n V_low
+ 792.300001n V_low
+ 792.400000n V_low
+ 792.400001n V_low
+ 792.500000n V_low
+ 792.500001n V_low
+ 792.600000n V_low
+ 792.600001n V_low
+ 792.700000n V_low
+ 792.700001n V_low
+ 792.800000n V_low
+ 792.800001n V_low
+ 792.900000n V_low
+ 792.900001n V_low
+ 793.000000n V_low
+ 793.000001n V_hig
+ 793.100000n V_hig
+ 793.100001n V_hig
+ 793.200000n V_hig
+ 793.200001n V_hig
+ 793.300000n V_hig
+ 793.300001n V_hig
+ 793.400000n V_hig
+ 793.400001n V_hig
+ 793.500000n V_hig
+ 793.500001n V_hig
+ 793.600000n V_hig
+ 793.600001n V_hig
+ 793.700000n V_hig
+ 793.700001n V_hig
+ 793.800000n V_hig
+ 793.800001n V_hig
+ 793.900000n V_hig
+ 793.900001n V_hig
+ 794.000000n V_hig
+ 794.000001n V_low
+ 794.100000n V_low
+ 794.100001n V_low
+ 794.200000n V_low
+ 794.200001n V_low
+ 794.300000n V_low
+ 794.300001n V_low
+ 794.400000n V_low
+ 794.400001n V_low
+ 794.500000n V_low
+ 794.500001n V_low
+ 794.600000n V_low
+ 794.600001n V_low
+ 794.700000n V_low
+ 794.700001n V_low
+ 794.800000n V_low
+ 794.800001n V_low
+ 794.900000n V_low
+ 794.900001n V_low
+ 795.000000n V_low
+ 795.000001n V_low
+ 795.100000n V_low
+ 795.100001n V_low
+ 795.200000n V_low
+ 795.200001n V_low
+ 795.300000n V_low
+ 795.300001n V_low
+ 795.400000n V_low
+ 795.400001n V_low
+ 795.500000n V_low
+ 795.500001n V_low
+ 795.600000n V_low
+ 795.600001n V_low
+ 795.700000n V_low
+ 795.700001n V_low
+ 795.800000n V_low
+ 795.800001n V_low
+ 795.900000n V_low
+ 795.900001n V_low
+ 796.000000n V_low
+ 796.000001n V_low
+ 796.100000n V_low
+ 796.100001n V_low
+ 796.200000n V_low
+ 796.200001n V_low
+ 796.300000n V_low
+ 796.300001n V_low
+ 796.400000n V_low
+ 796.400001n V_low
+ 796.500000n V_low
+ 796.500001n V_low
+ 796.600000n V_low
+ 796.600001n V_low
+ 796.700000n V_low
+ 796.700001n V_low
+ 796.800000n V_low
+ 796.800001n V_low
+ 796.900000n V_low
+ 796.900001n V_low
+ 797.000000n V_low
+ 797.000001n V_low
+ 797.100000n V_low
+ 797.100001n V_low
+ 797.200000n V_low
+ 797.200001n V_low
+ 797.300000n V_low
+ 797.300001n V_low
+ 797.400000n V_low
+ 797.400001n V_low
+ 797.500000n V_low
+ 797.500001n V_low
+ 797.600000n V_low
+ 797.600001n V_low
+ 797.700000n V_low
+ 797.700001n V_low
+ 797.800000n V_low
+ 797.800001n V_low
+ 797.900000n V_low
+ 797.900001n V_low
+ 798.000000n V_low
+ 798.000001n V_hig
+ 798.100000n V_hig
+ 798.100001n V_hig
+ 798.200000n V_hig
+ 798.200001n V_hig
+ 798.300000n V_hig
+ 798.300001n V_hig
+ 798.400000n V_hig
+ 798.400001n V_hig
+ 798.500000n V_hig
+ 798.500001n V_hig
+ 798.600000n V_hig
+ 798.600001n V_hig
+ 798.700000n V_hig
+ 798.700001n V_hig
+ 798.800000n V_hig
+ 798.800001n V_hig
+ 798.900000n V_hig
+ 798.900001n V_hig
+ 799.000000n V_hig
+ 799.000001n V_low
+ 799.100000n V_low
+ 799.100001n V_low
+ 799.200000n V_low
+ 799.200001n V_low
+ 799.300000n V_low
+ 799.300001n V_low
+ 799.400000n V_low
+ 799.400001n V_low
+ 799.500000n V_low
+ 799.500001n V_low
+ 799.600000n V_low
+ 799.600001n V_low
+ 799.700000n V_low
+ 799.700001n V_low
+ 799.800000n V_low
+ 799.800001n V_low
+ 799.900000n V_low
+ 799.900001n V_low
+ 800.000000n V_low
+ 800.000001n V_hig
+ 800.100000n V_hig
+ 800.100001n V_hig
+ 800.200000n V_hig
+ 800.200001n V_hig
+ 800.300000n V_hig
+ 800.300001n V_hig
+ 800.400000n V_hig
+ 800.400001n V_hig
+ 800.500000n V_hig
+ 800.500001n V_hig
+ 800.600000n V_hig
+ 800.600001n V_hig
+ 800.700000n V_hig
+ 800.700001n V_hig
+ 800.800000n V_hig
+ 800.800001n V_hig
+ 800.900000n V_hig
+ 800.900001n V_hig
+ 801.000000n V_hig
+ 801.000001n V_low
+ 801.100000n V_low
+ 801.100001n V_low
+ 801.200000n V_low
+ 801.200001n V_low
+ 801.300000n V_low
+ 801.300001n V_low
+ 801.400000n V_low
+ 801.400001n V_low
+ 801.500000n V_low
+ 801.500001n V_low
+ 801.600000n V_low
+ 801.600001n V_low
+ 801.700000n V_low
+ 801.700001n V_low
+ 801.800000n V_low
+ 801.800001n V_low
+ 801.900000n V_low
+ 801.900001n V_low
+ 802.000000n V_low
+ 802.000001n V_low
+ 802.100000n V_low
+ 802.100001n V_low
+ 802.200000n V_low
+ 802.200001n V_low
+ 802.300000n V_low
+ 802.300001n V_low
+ 802.400000n V_low
+ 802.400001n V_low
+ 802.500000n V_low
+ 802.500001n V_low
+ 802.600000n V_low
+ 802.600001n V_low
+ 802.700000n V_low
+ 802.700001n V_low
+ 802.800000n V_low
+ 802.800001n V_low
+ 802.900000n V_low
+ 802.900001n V_low
+ 803.000000n V_low
+ 803.000001n V_low
+ 803.100000n V_low
+ 803.100001n V_low
+ 803.200000n V_low
+ 803.200001n V_low
+ 803.300000n V_low
+ 803.300001n V_low
+ 803.400000n V_low
+ 803.400001n V_low
+ 803.500000n V_low
+ 803.500001n V_low
+ 803.600000n V_low
+ 803.600001n V_low
+ 803.700000n V_low
+ 803.700001n V_low
+ 803.800000n V_low
+ 803.800001n V_low
+ 803.900000n V_low
+ 803.900001n V_low
+ 804.000000n V_low
+ 804.000001n V_low
+ 804.100000n V_low
+ 804.100001n V_low
+ 804.200000n V_low
+ 804.200001n V_low
+ 804.300000n V_low
+ 804.300001n V_low
+ 804.400000n V_low
+ 804.400001n V_low
+ 804.500000n V_low
+ 804.500001n V_low
+ 804.600000n V_low
+ 804.600001n V_low
+ 804.700000n V_low
+ 804.700001n V_low
+ 804.800000n V_low
+ 804.800001n V_low
+ 804.900000n V_low
+ 804.900001n V_low
+ 805.000000n V_low
+ 805.000001n V_low
+ 805.100000n V_low
+ 805.100001n V_low
+ 805.200000n V_low
+ 805.200001n V_low
+ 805.300000n V_low
+ 805.300001n V_low
+ 805.400000n V_low
+ 805.400001n V_low
+ 805.500000n V_low
+ 805.500001n V_low
+ 805.600000n V_low
+ 805.600001n V_low
+ 805.700000n V_low
+ 805.700001n V_low
+ 805.800000n V_low
+ 805.800001n V_low
+ 805.900000n V_low
+ 805.900001n V_low
+ 806.000000n V_low
+ 806.000001n V_hig
+ 806.100000n V_hig
+ 806.100001n V_hig
+ 806.200000n V_hig
+ 806.200001n V_hig
+ 806.300000n V_hig
+ 806.300001n V_hig
+ 806.400000n V_hig
+ 806.400001n V_hig
+ 806.500000n V_hig
+ 806.500001n V_hig
+ 806.600000n V_hig
+ 806.600001n V_hig
+ 806.700000n V_hig
+ 806.700001n V_hig
+ 806.800000n V_hig
+ 806.800001n V_hig
+ 806.900000n V_hig
+ 806.900001n V_hig
+ 807.000000n V_hig
+ 807.000001n V_low
+ 807.100000n V_low
+ 807.100001n V_low
+ 807.200000n V_low
+ 807.200001n V_low
+ 807.300000n V_low
+ 807.300001n V_low
+ 807.400000n V_low
+ 807.400001n V_low
+ 807.500000n V_low
+ 807.500001n V_low
+ 807.600000n V_low
+ 807.600001n V_low
+ 807.700000n V_low
+ 807.700001n V_low
+ 807.800000n V_low
+ 807.800001n V_low
+ 807.900000n V_low
+ 807.900001n V_low
+ 808.000000n V_low
+ 808.000001n V_hig
+ 808.100000n V_hig
+ 808.100001n V_hig
+ 808.200000n V_hig
+ 808.200001n V_hig
+ 808.300000n V_hig
+ 808.300001n V_hig
+ 808.400000n V_hig
+ 808.400001n V_hig
+ 808.500000n V_hig
+ 808.500001n V_hig
+ 808.600000n V_hig
+ 808.600001n V_hig
+ 808.700000n V_hig
+ 808.700001n V_hig
+ 808.800000n V_hig
+ 808.800001n V_hig
+ 808.900000n V_hig
+ 808.900001n V_hig
+ 809.000000n V_hig
+ 809.000001n V_hig
+ 809.100000n V_hig
+ 809.100001n V_hig
+ 809.200000n V_hig
+ 809.200001n V_hig
+ 809.300000n V_hig
+ 809.300001n V_hig
+ 809.400000n V_hig
+ 809.400001n V_hig
+ 809.500000n V_hig
+ 809.500001n V_hig
+ 809.600000n V_hig
+ 809.600001n V_hig
+ 809.700000n V_hig
+ 809.700001n V_hig
+ 809.800000n V_hig
+ 809.800001n V_hig
+ 809.900000n V_hig
+ 809.900001n V_hig
+ 810.000000n V_hig
+ 810.000001n V_low
+ 810.100000n V_low
+ 810.100001n V_low
+ 810.200000n V_low
+ 810.200001n V_low
+ 810.300000n V_low
+ 810.300001n V_low
+ 810.400000n V_low
+ 810.400001n V_low
+ 810.500000n V_low
+ 810.500001n V_low
+ 810.600000n V_low
+ 810.600001n V_low
+ 810.700000n V_low
+ 810.700001n V_low
+ 810.800000n V_low
+ 810.800001n V_low
+ 810.900000n V_low
+ 810.900001n V_low
+ 811.000000n V_low
+ 811.000001n V_hig
+ 811.100000n V_hig
+ 811.100001n V_hig
+ 811.200000n V_hig
+ 811.200001n V_hig
+ 811.300000n V_hig
+ 811.300001n V_hig
+ 811.400000n V_hig
+ 811.400001n V_hig
+ 811.500000n V_hig
+ 811.500001n V_hig
+ 811.600000n V_hig
+ 811.600001n V_hig
+ 811.700000n V_hig
+ 811.700001n V_hig
+ 811.800000n V_hig
+ 811.800001n V_hig
+ 811.900000n V_hig
+ 811.900001n V_hig
+ 812.000000n V_hig
+ 812.000001n V_low
+ 812.100000n V_low
+ 812.100001n V_low
+ 812.200000n V_low
+ 812.200001n V_low
+ 812.300000n V_low
+ 812.300001n V_low
+ 812.400000n V_low
+ 812.400001n V_low
+ 812.500000n V_low
+ 812.500001n V_low
+ 812.600000n V_low
+ 812.600001n V_low
+ 812.700000n V_low
+ 812.700001n V_low
+ 812.800000n V_low
+ 812.800001n V_low
+ 812.900000n V_low
+ 812.900001n V_low
+ 813.000000n V_low
+ 813.000001n V_hig
+ 813.100000n V_hig
+ 813.100001n V_hig
+ 813.200000n V_hig
+ 813.200001n V_hig
+ 813.300000n V_hig
+ 813.300001n V_hig
+ 813.400000n V_hig
+ 813.400001n V_hig
+ 813.500000n V_hig
+ 813.500001n V_hig
+ 813.600000n V_hig
+ 813.600001n V_hig
+ 813.700000n V_hig
+ 813.700001n V_hig
+ 813.800000n V_hig
+ 813.800001n V_hig
+ 813.900000n V_hig
+ 813.900001n V_hig
+ 814.000000n V_hig
+ 814.000001n V_low
+ 814.100000n V_low
+ 814.100001n V_low
+ 814.200000n V_low
+ 814.200001n V_low
+ 814.300000n V_low
+ 814.300001n V_low
+ 814.400000n V_low
+ 814.400001n V_low
+ 814.500000n V_low
+ 814.500001n V_low
+ 814.600000n V_low
+ 814.600001n V_low
+ 814.700000n V_low
+ 814.700001n V_low
+ 814.800000n V_low
+ 814.800001n V_low
+ 814.900000n V_low
+ 814.900001n V_low
+ 815.000000n V_low
+ 815.000001n V_low
+ 815.100000n V_low
+ 815.100001n V_low
+ 815.200000n V_low
+ 815.200001n V_low
+ 815.300000n V_low
+ 815.300001n V_low
+ 815.400000n V_low
+ 815.400001n V_low
+ 815.500000n V_low
+ 815.500001n V_low
+ 815.600000n V_low
+ 815.600001n V_low
+ 815.700000n V_low
+ 815.700001n V_low
+ 815.800000n V_low
+ 815.800001n V_low
+ 815.900000n V_low
+ 815.900001n V_low
+ 816.000000n V_low
+ 816.000001n V_low
+ 816.100000n V_low
+ 816.100001n V_low
+ 816.200000n V_low
+ 816.200001n V_low
+ 816.300000n V_low
+ 816.300001n V_low
+ 816.400000n V_low
+ 816.400001n V_low
+ 816.500000n V_low
+ 816.500001n V_low
+ 816.600000n V_low
+ 816.600001n V_low
+ 816.700000n V_low
+ 816.700001n V_low
+ 816.800000n V_low
+ 816.800001n V_low
+ 816.900000n V_low
+ 816.900001n V_low
+ 817.000000n V_low
+ 817.000001n V_hig
+ 817.100000n V_hig
+ 817.100001n V_hig
+ 817.200000n V_hig
+ 817.200001n V_hig
+ 817.300000n V_hig
+ 817.300001n V_hig
+ 817.400000n V_hig
+ 817.400001n V_hig
+ 817.500000n V_hig
+ 817.500001n V_hig
+ 817.600000n V_hig
+ 817.600001n V_hig
+ 817.700000n V_hig
+ 817.700001n V_hig
+ 817.800000n V_hig
+ 817.800001n V_hig
+ 817.900000n V_hig
+ 817.900001n V_hig
+ 818.000000n V_hig
+ 818.000001n V_low
+ 818.100000n V_low
+ 818.100001n V_low
+ 818.200000n V_low
+ 818.200001n V_low
+ 818.300000n V_low
+ 818.300001n V_low
+ 818.400000n V_low
+ 818.400001n V_low
+ 818.500000n V_low
+ 818.500001n V_low
+ 818.600000n V_low
+ 818.600001n V_low
+ 818.700000n V_low
+ 818.700001n V_low
+ 818.800000n V_low
+ 818.800001n V_low
+ 818.900000n V_low
+ 818.900001n V_low
+ 819.000000n V_low
+ 819.000001n V_low
+ 819.100000n V_low
+ 819.100001n V_low
+ 819.200000n V_low
+ 819.200001n V_low
+ 819.300000n V_low
+ 819.300001n V_low
+ 819.400000n V_low
+ 819.400001n V_low
+ 819.500000n V_low
+ 819.500001n V_low
+ 819.600000n V_low
+ 819.600001n V_low
+ 819.700000n V_low
+ 819.700001n V_low
+ 819.800000n V_low
+ 819.800001n V_low
+ 819.900000n V_low
+ 819.900001n V_low
+ 820.000000n V_low
+ 820.000001n V_low
+ 820.100000n V_low
+ 820.100001n V_low
+ 820.200000n V_low
+ 820.200001n V_low
+ 820.300000n V_low
+ 820.300001n V_low
+ 820.400000n V_low
+ 820.400001n V_low
+ 820.500000n V_low
+ 820.500001n V_low
+ 820.600000n V_low
+ 820.600001n V_low
+ 820.700000n V_low
+ 820.700001n V_low
+ 820.800000n V_low
+ 820.800001n V_low
+ 820.900000n V_low
+ 820.900001n V_low
+ 821.000000n V_low
+ 821.000001n V_hig
+ 821.100000n V_hig
+ 821.100001n V_hig
+ 821.200000n V_hig
+ 821.200001n V_hig
+ 821.300000n V_hig
+ 821.300001n V_hig
+ 821.400000n V_hig
+ 821.400001n V_hig
+ 821.500000n V_hig
+ 821.500001n V_hig
+ 821.600000n V_hig
+ 821.600001n V_hig
+ 821.700000n V_hig
+ 821.700001n V_hig
+ 821.800000n V_hig
+ 821.800001n V_hig
+ 821.900000n V_hig
+ 821.900001n V_hig
+ 822.000000n V_hig
+ 822.000001n V_low
+ 822.100000n V_low
+ 822.100001n V_low
+ 822.200000n V_low
+ 822.200001n V_low
+ 822.300000n V_low
+ 822.300001n V_low
+ 822.400000n V_low
+ 822.400001n V_low
+ 822.500000n V_low
+ 822.500001n V_low
+ 822.600000n V_low
+ 822.600001n V_low
+ 822.700000n V_low
+ 822.700001n V_low
+ 822.800000n V_low
+ 822.800001n V_low
+ 822.900000n V_low
+ 822.900001n V_low
+ 823.000000n V_low
+ 823.000001n V_low
+ 823.100000n V_low
+ 823.100001n V_low
+ 823.200000n V_low
+ 823.200001n V_low
+ 823.300000n V_low
+ 823.300001n V_low
+ 823.400000n V_low
+ 823.400001n V_low
+ 823.500000n V_low
+ 823.500001n V_low
+ 823.600000n V_low
+ 823.600001n V_low
+ 823.700000n V_low
+ 823.700001n V_low
+ 823.800000n V_low
+ 823.800001n V_low
+ 823.900000n V_low
+ 823.900001n V_low
+ 824.000000n V_low
+ 824.000001n V_hig
+ 824.100000n V_hig
+ 824.100001n V_hig
+ 824.200000n V_hig
+ 824.200001n V_hig
+ 824.300000n V_hig
+ 824.300001n V_hig
+ 824.400000n V_hig
+ 824.400001n V_hig
+ 824.500000n V_hig
+ 824.500001n V_hig
+ 824.600000n V_hig
+ 824.600001n V_hig
+ 824.700000n V_hig
+ 824.700001n V_hig
+ 824.800000n V_hig
+ 824.800001n V_hig
+ 824.900000n V_hig
+ 824.900001n V_hig
+ 825.000000n V_hig
+ 825.000001n V_low
+ 825.100000n V_low
+ 825.100001n V_low
+ 825.200000n V_low
+ 825.200001n V_low
+ 825.300000n V_low
+ 825.300001n V_low
+ 825.400000n V_low
+ 825.400001n V_low
+ 825.500000n V_low
+ 825.500001n V_low
+ 825.600000n V_low
+ 825.600001n V_low
+ 825.700000n V_low
+ 825.700001n V_low
+ 825.800000n V_low
+ 825.800001n V_low
+ 825.900000n V_low
+ 825.900001n V_low
+ 826.000000n V_low
+ 826.000001n V_hig
+ 826.100000n V_hig
+ 826.100001n V_hig
+ 826.200000n V_hig
+ 826.200001n V_hig
+ 826.300000n V_hig
+ 826.300001n V_hig
+ 826.400000n V_hig
+ 826.400001n V_hig
+ 826.500000n V_hig
+ 826.500001n V_hig
+ 826.600000n V_hig
+ 826.600001n V_hig
+ 826.700000n V_hig
+ 826.700001n V_hig
+ 826.800000n V_hig
+ 826.800001n V_hig
+ 826.900000n V_hig
+ 826.900001n V_hig
+ 827.000000n V_hig
+ 827.000001n V_hig
+ 827.100000n V_hig
+ 827.100001n V_hig
+ 827.200000n V_hig
+ 827.200001n V_hig
+ 827.300000n V_hig
+ 827.300001n V_hig
+ 827.400000n V_hig
+ 827.400001n V_hig
+ 827.500000n V_hig
+ 827.500001n V_hig
+ 827.600000n V_hig
+ 827.600001n V_hig
+ 827.700000n V_hig
+ 827.700001n V_hig
+ 827.800000n V_hig
+ 827.800001n V_hig
+ 827.900000n V_hig
+ 827.900001n V_hig
+ 828.000000n V_hig
+ 828.000001n V_low
+ 828.100000n V_low
+ 828.100001n V_low
+ 828.200000n V_low
+ 828.200001n V_low
+ 828.300000n V_low
+ 828.300001n V_low
+ 828.400000n V_low
+ 828.400001n V_low
+ 828.500000n V_low
+ 828.500001n V_low
+ 828.600000n V_low
+ 828.600001n V_low
+ 828.700000n V_low
+ 828.700001n V_low
+ 828.800000n V_low
+ 828.800001n V_low
+ 828.900000n V_low
+ 828.900001n V_low
+ 829.000000n V_low
+ 829.000001n V_low
+ 829.100000n V_low
+ 829.100001n V_low
+ 829.200000n V_low
+ 829.200001n V_low
+ 829.300000n V_low
+ 829.300001n V_low
+ 829.400000n V_low
+ 829.400001n V_low
+ 829.500000n V_low
+ 829.500001n V_low
+ 829.600000n V_low
+ 829.600001n V_low
+ 829.700000n V_low
+ 829.700001n V_low
+ 829.800000n V_low
+ 829.800001n V_low
+ 829.900000n V_low
+ 829.900001n V_low
+ 830.000000n V_low
+ 830.000001n V_low
+ 830.100000n V_low
+ 830.100001n V_low
+ 830.200000n V_low
+ 830.200001n V_low
+ 830.300000n V_low
+ 830.300001n V_low
+ 830.400000n V_low
+ 830.400001n V_low
+ 830.500000n V_low
+ 830.500001n V_low
+ 830.600000n V_low
+ 830.600001n V_low
+ 830.700000n V_low
+ 830.700001n V_low
+ 830.800000n V_low
+ 830.800001n V_low
+ 830.900000n V_low
+ 830.900001n V_low
+ 831.000000n V_low
+ 831.000001n V_low
+ 831.100000n V_low
+ 831.100001n V_low
+ 831.200000n V_low
+ 831.200001n V_low
+ 831.300000n V_low
+ 831.300001n V_low
+ 831.400000n V_low
+ 831.400001n V_low
+ 831.500000n V_low
+ 831.500001n V_low
+ 831.600000n V_low
+ 831.600001n V_low
+ 831.700000n V_low
+ 831.700001n V_low
+ 831.800000n V_low
+ 831.800001n V_low
+ 831.900000n V_low
+ 831.900001n V_low
+ 832.000000n V_low
+ 832.000001n V_hig
+ 832.100000n V_hig
+ 832.100001n V_hig
+ 832.200000n V_hig
+ 832.200001n V_hig
+ 832.300000n V_hig
+ 832.300001n V_hig
+ 832.400000n V_hig
+ 832.400001n V_hig
+ 832.500000n V_hig
+ 832.500001n V_hig
+ 832.600000n V_hig
+ 832.600001n V_hig
+ 832.700000n V_hig
+ 832.700001n V_hig
+ 832.800000n V_hig
+ 832.800001n V_hig
+ 832.900000n V_hig
+ 832.900001n V_hig
+ 833.000000n V_hig
+ 833.000001n V_hig
+ 833.100000n V_hig
+ 833.100001n V_hig
+ 833.200000n V_hig
+ 833.200001n V_hig
+ 833.300000n V_hig
+ 833.300001n V_hig
+ 833.400000n V_hig
+ 833.400001n V_hig
+ 833.500000n V_hig
+ 833.500001n V_hig
+ 833.600000n V_hig
+ 833.600001n V_hig
+ 833.700000n V_hig
+ 833.700001n V_hig
+ 833.800000n V_hig
+ 833.800001n V_hig
+ 833.900000n V_hig
+ 833.900001n V_hig
+ 834.000000n V_hig
+ 834.000001n V_low
+ 834.100000n V_low
+ 834.100001n V_low
+ 834.200000n V_low
+ 834.200001n V_low
+ 834.300000n V_low
+ 834.300001n V_low
+ 834.400000n V_low
+ 834.400001n V_low
+ 834.500000n V_low
+ 834.500001n V_low
+ 834.600000n V_low
+ 834.600001n V_low
+ 834.700000n V_low
+ 834.700001n V_low
+ 834.800000n V_low
+ 834.800001n V_low
+ 834.900000n V_low
+ 834.900001n V_low
+ 835.000000n V_low
+ 835.000001n V_low
+ 835.100000n V_low
+ 835.100001n V_low
+ 835.200000n V_low
+ 835.200001n V_low
+ 835.300000n V_low
+ 835.300001n V_low
+ 835.400000n V_low
+ 835.400001n V_low
+ 835.500000n V_low
+ 835.500001n V_low
+ 835.600000n V_low
+ 835.600001n V_low
+ 835.700000n V_low
+ 835.700001n V_low
+ 835.800000n V_low
+ 835.800001n V_low
+ 835.900000n V_low
+ 835.900001n V_low
+ 836.000000n V_low
+ 836.000001n V_low
+ 836.100000n V_low
+ 836.100001n V_low
+ 836.200000n V_low
+ 836.200001n V_low
+ 836.300000n V_low
+ 836.300001n V_low
+ 836.400000n V_low
+ 836.400001n V_low
+ 836.500000n V_low
+ 836.500001n V_low
+ 836.600000n V_low
+ 836.600001n V_low
+ 836.700000n V_low
+ 836.700001n V_low
+ 836.800000n V_low
+ 836.800001n V_low
+ 836.900000n V_low
+ 836.900001n V_low
+ 837.000000n V_low
+ 837.000001n V_low
+ 837.100000n V_low
+ 837.100001n V_low
+ 837.200000n V_low
+ 837.200001n V_low
+ 837.300000n V_low
+ 837.300001n V_low
+ 837.400000n V_low
+ 837.400001n V_low
+ 837.500000n V_low
+ 837.500001n V_low
+ 837.600000n V_low
+ 837.600001n V_low
+ 837.700000n V_low
+ 837.700001n V_low
+ 837.800000n V_low
+ 837.800001n V_low
+ 837.900000n V_low
+ 837.900001n V_low
+ 838.000000n V_low
+ 838.000001n V_hig
+ 838.100000n V_hig
+ 838.100001n V_hig
+ 838.200000n V_hig
+ 838.200001n V_hig
+ 838.300000n V_hig
+ 838.300001n V_hig
+ 838.400000n V_hig
+ 838.400001n V_hig
+ 838.500000n V_hig
+ 838.500001n V_hig
+ 838.600000n V_hig
+ 838.600001n V_hig
+ 838.700000n V_hig
+ 838.700001n V_hig
+ 838.800000n V_hig
+ 838.800001n V_hig
+ 838.900000n V_hig
+ 838.900001n V_hig
+ 839.000000n V_hig
+ 839.000001n V_hig
+ 839.100000n V_hig
+ 839.100001n V_hig
+ 839.200000n V_hig
+ 839.200001n V_hig
+ 839.300000n V_hig
+ 839.300001n V_hig
+ 839.400000n V_hig
+ 839.400001n V_hig
+ 839.500000n V_hig
+ 839.500001n V_hig
+ 839.600000n V_hig
+ 839.600001n V_hig
+ 839.700000n V_hig
+ 839.700001n V_hig
+ 839.800000n V_hig
+ 839.800001n V_hig
+ 839.900000n V_hig
+ 839.900001n V_hig
+ 840.000000n V_hig
+ 840.000001n V_low
+ 840.100000n V_low
+ 840.100001n V_low
+ 840.200000n V_low
+ 840.200001n V_low
+ 840.300000n V_low
+ 840.300001n V_low
+ 840.400000n V_low
+ 840.400001n V_low
+ 840.500000n V_low
+ 840.500001n V_low
+ 840.600000n V_low
+ 840.600001n V_low
+ 840.700000n V_low
+ 840.700001n V_low
+ 840.800000n V_low
+ 840.800001n V_low
+ 840.900000n V_low
+ 840.900001n V_low
+ 841.000000n V_low
+ 841.000001n V_hig
+ 841.100000n V_hig
+ 841.100001n V_hig
+ 841.200000n V_hig
+ 841.200001n V_hig
+ 841.300000n V_hig
+ 841.300001n V_hig
+ 841.400000n V_hig
+ 841.400001n V_hig
+ 841.500000n V_hig
+ 841.500001n V_hig
+ 841.600000n V_hig
+ 841.600001n V_hig
+ 841.700000n V_hig
+ 841.700001n V_hig
+ 841.800000n V_hig
+ 841.800001n V_hig
+ 841.900000n V_hig
+ 841.900001n V_hig
+ 842.000000n V_hig
+ 842.000001n V_hig
+ 842.100000n V_hig
+ 842.100001n V_hig
+ 842.200000n V_hig
+ 842.200001n V_hig
+ 842.300000n V_hig
+ 842.300001n V_hig
+ 842.400000n V_hig
+ 842.400001n V_hig
+ 842.500000n V_hig
+ 842.500001n V_hig
+ 842.600000n V_hig
+ 842.600001n V_hig
+ 842.700000n V_hig
+ 842.700001n V_hig
+ 842.800000n V_hig
+ 842.800001n V_hig
+ 842.900000n V_hig
+ 842.900001n V_hig
+ 843.000000n V_hig
+ 843.000001n V_hig
+ 843.100000n V_hig
+ 843.100001n V_hig
+ 843.200000n V_hig
+ 843.200001n V_hig
+ 843.300000n V_hig
+ 843.300001n V_hig
+ 843.400000n V_hig
+ 843.400001n V_hig
+ 843.500000n V_hig
+ 843.500001n V_hig
+ 843.600000n V_hig
+ 843.600001n V_hig
+ 843.700000n V_hig
+ 843.700001n V_hig
+ 843.800000n V_hig
+ 843.800001n V_hig
+ 843.900000n V_hig
+ 843.900001n V_hig
+ 844.000000n V_hig
+ 844.000001n V_hig
+ 844.100000n V_hig
+ 844.100001n V_hig
+ 844.200000n V_hig
+ 844.200001n V_hig
+ 844.300000n V_hig
+ 844.300001n V_hig
+ 844.400000n V_hig
+ 844.400001n V_hig
+ 844.500000n V_hig
+ 844.500001n V_hig
+ 844.600000n V_hig
+ 844.600001n V_hig
+ 844.700000n V_hig
+ 844.700001n V_hig
+ 844.800000n V_hig
+ 844.800001n V_hig
+ 844.900000n V_hig
+ 844.900001n V_hig
+ 845.000000n V_hig
+ 845.000001n V_hig
+ 845.100000n V_hig
+ 845.100001n V_hig
+ 845.200000n V_hig
+ 845.200001n V_hig
+ 845.300000n V_hig
+ 845.300001n V_hig
+ 845.400000n V_hig
+ 845.400001n V_hig
+ 845.500000n V_hig
+ 845.500001n V_hig
+ 845.600000n V_hig
+ 845.600001n V_hig
+ 845.700000n V_hig
+ 845.700001n V_hig
+ 845.800000n V_hig
+ 845.800001n V_hig
+ 845.900000n V_hig
+ 845.900001n V_hig
+ 846.000000n V_hig
+ 846.000001n V_low
+ 846.100000n V_low
+ 846.100001n V_low
+ 846.200000n V_low
+ 846.200001n V_low
+ 846.300000n V_low
+ 846.300001n V_low
+ 846.400000n V_low
+ 846.400001n V_low
+ 846.500000n V_low
+ 846.500001n V_low
+ 846.600000n V_low
+ 846.600001n V_low
+ 846.700000n V_low
+ 846.700001n V_low
+ 846.800000n V_low
+ 846.800001n V_low
+ 846.900000n V_low
+ 846.900001n V_low
+ 847.000000n V_low
+ 847.000001n V_hig
+ 847.100000n V_hig
+ 847.100001n V_hig
+ 847.200000n V_hig
+ 847.200001n V_hig
+ 847.300000n V_hig
+ 847.300001n V_hig
+ 847.400000n V_hig
+ 847.400001n V_hig
+ 847.500000n V_hig
+ 847.500001n V_hig
+ 847.600000n V_hig
+ 847.600001n V_hig
+ 847.700000n V_hig
+ 847.700001n V_hig
+ 847.800000n V_hig
+ 847.800001n V_hig
+ 847.900000n V_hig
+ 847.900001n V_hig
+ 848.000000n V_hig
+ 848.000001n V_hig
+ 848.100000n V_hig
+ 848.100001n V_hig
+ 848.200000n V_hig
+ 848.200001n V_hig
+ 848.300000n V_hig
+ 848.300001n V_hig
+ 848.400000n V_hig
+ 848.400001n V_hig
+ 848.500000n V_hig
+ 848.500001n V_hig
+ 848.600000n V_hig
+ 848.600001n V_hig
+ 848.700000n V_hig
+ 848.700001n V_hig
+ 848.800000n V_hig
+ 848.800001n V_hig
+ 848.900000n V_hig
+ 848.900001n V_hig
+ 849.000000n V_hig
+ 849.000001n V_hig
+ 849.100000n V_hig
+ 849.100001n V_hig
+ 849.200000n V_hig
+ 849.200001n V_hig
+ 849.300000n V_hig
+ 849.300001n V_hig
+ 849.400000n V_hig
+ 849.400001n V_hig
+ 849.500000n V_hig
+ 849.500001n V_hig
+ 849.600000n V_hig
+ 849.600001n V_hig
+ 849.700000n V_hig
+ 849.700001n V_hig
+ 849.800000n V_hig
+ 849.800001n V_hig
+ 849.900000n V_hig
+ 849.900001n V_hig
+ 850.000000n V_hig
+ 850.000001n V_hig
+ 850.100000n V_hig
+ 850.100001n V_hig
+ 850.200000n V_hig
+ 850.200001n V_hig
+ 850.300000n V_hig
+ 850.300001n V_hig
+ 850.400000n V_hig
+ 850.400001n V_hig
+ 850.500000n V_hig
+ 850.500001n V_hig
+ 850.600000n V_hig
+ 850.600001n V_hig
+ 850.700000n V_hig
+ 850.700001n V_hig
+ 850.800000n V_hig
+ 850.800001n V_hig
+ 850.900000n V_hig
+ 850.900001n V_hig
+ 851.000000n V_hig
+ 851.000001n V_hig
+ 851.100000n V_hig
+ 851.100001n V_hig
+ 851.200000n V_hig
+ 851.200001n V_hig
+ 851.300000n V_hig
+ 851.300001n V_hig
+ 851.400000n V_hig
+ 851.400001n V_hig
+ 851.500000n V_hig
+ 851.500001n V_hig
+ 851.600000n V_hig
+ 851.600001n V_hig
+ 851.700000n V_hig
+ 851.700001n V_hig
+ 851.800000n V_hig
+ 851.800001n V_hig
+ 851.900000n V_hig
+ 851.900001n V_hig
+ 852.000000n V_hig
+ 852.000001n V_low
+ 852.100000n V_low
+ 852.100001n V_low
+ 852.200000n V_low
+ 852.200001n V_low
+ 852.300000n V_low
+ 852.300001n V_low
+ 852.400000n V_low
+ 852.400001n V_low
+ 852.500000n V_low
+ 852.500001n V_low
+ 852.600000n V_low
+ 852.600001n V_low
+ 852.700000n V_low
+ 852.700001n V_low
+ 852.800000n V_low
+ 852.800001n V_low
+ 852.900000n V_low
+ 852.900001n V_low
+ 853.000000n V_low
+ 853.000001n V_hig
+ 853.100000n V_hig
+ 853.100001n V_hig
+ 853.200000n V_hig
+ 853.200001n V_hig
+ 853.300000n V_hig
+ 853.300001n V_hig
+ 853.400000n V_hig
+ 853.400001n V_hig
+ 853.500000n V_hig
+ 853.500001n V_hig
+ 853.600000n V_hig
+ 853.600001n V_hig
+ 853.700000n V_hig
+ 853.700001n V_hig
+ 853.800000n V_hig
+ 853.800001n V_hig
+ 853.900000n V_hig
+ 853.900001n V_hig
+ 854.000000n V_hig
+ 854.000001n V_hig
+ 854.100000n V_hig
+ 854.100001n V_hig
+ 854.200000n V_hig
+ 854.200001n V_hig
+ 854.300000n V_hig
+ 854.300001n V_hig
+ 854.400000n V_hig
+ 854.400001n V_hig
+ 854.500000n V_hig
+ 854.500001n V_hig
+ 854.600000n V_hig
+ 854.600001n V_hig
+ 854.700000n V_hig
+ 854.700001n V_hig
+ 854.800000n V_hig
+ 854.800001n V_hig
+ 854.900000n V_hig
+ 854.900001n V_hig
+ 855.000000n V_hig
+ 855.000001n V_hig
+ 855.100000n V_hig
+ 855.100001n V_hig
+ 855.200000n V_hig
+ 855.200001n V_hig
+ 855.300000n V_hig
+ 855.300001n V_hig
+ 855.400000n V_hig
+ 855.400001n V_hig
+ 855.500000n V_hig
+ 855.500001n V_hig
+ 855.600000n V_hig
+ 855.600001n V_hig
+ 855.700000n V_hig
+ 855.700001n V_hig
+ 855.800000n V_hig
+ 855.800001n V_hig
+ 855.900000n V_hig
+ 855.900001n V_hig
+ 856.000000n V_hig
+ 856.000001n V_low
+ 856.100000n V_low
+ 856.100001n V_low
+ 856.200000n V_low
+ 856.200001n V_low
+ 856.300000n V_low
+ 856.300001n V_low
+ 856.400000n V_low
+ 856.400001n V_low
+ 856.500000n V_low
+ 856.500001n V_low
+ 856.600000n V_low
+ 856.600001n V_low
+ 856.700000n V_low
+ 856.700001n V_low
+ 856.800000n V_low
+ 856.800001n V_low
+ 856.900000n V_low
+ 856.900001n V_low
+ 857.000000n V_low
+ 857.000001n V_hig
+ 857.100000n V_hig
+ 857.100001n V_hig
+ 857.200000n V_hig
+ 857.200001n V_hig
+ 857.300000n V_hig
+ 857.300001n V_hig
+ 857.400000n V_hig
+ 857.400001n V_hig
+ 857.500000n V_hig
+ 857.500001n V_hig
+ 857.600000n V_hig
+ 857.600001n V_hig
+ 857.700000n V_hig
+ 857.700001n V_hig
+ 857.800000n V_hig
+ 857.800001n V_hig
+ 857.900000n V_hig
+ 857.900001n V_hig
+ 858.000000n V_hig
+ 858.000001n V_low
+ 858.100000n V_low
+ 858.100001n V_low
+ 858.200000n V_low
+ 858.200001n V_low
+ 858.300000n V_low
+ 858.300001n V_low
+ 858.400000n V_low
+ 858.400001n V_low
+ 858.500000n V_low
+ 858.500001n V_low
+ 858.600000n V_low
+ 858.600001n V_low
+ 858.700000n V_low
+ 858.700001n V_low
+ 858.800000n V_low
+ 858.800001n V_low
+ 858.900000n V_low
+ 858.900001n V_low
+ 859.000000n V_low
+ 859.000001n V_hig
+ 859.100000n V_hig
+ 859.100001n V_hig
+ 859.200000n V_hig
+ 859.200001n V_hig
+ 859.300000n V_hig
+ 859.300001n V_hig
+ 859.400000n V_hig
+ 859.400001n V_hig
+ 859.500000n V_hig
+ 859.500001n V_hig
+ 859.600000n V_hig
+ 859.600001n V_hig
+ 859.700000n V_hig
+ 859.700001n V_hig
+ 859.800000n V_hig
+ 859.800001n V_hig
+ 859.900000n V_hig
+ 859.900001n V_hig
+ 860.000000n V_hig
+ 860.000001n V_low
+ 860.100000n V_low
+ 860.100001n V_low
+ 860.200000n V_low
+ 860.200001n V_low
+ 860.300000n V_low
+ 860.300001n V_low
+ 860.400000n V_low
+ 860.400001n V_low
+ 860.500000n V_low
+ 860.500001n V_low
+ 860.600000n V_low
+ 860.600001n V_low
+ 860.700000n V_low
+ 860.700001n V_low
+ 860.800000n V_low
+ 860.800001n V_low
+ 860.900000n V_low
+ 860.900001n V_low
+ 861.000000n V_low
+ 861.000001n V_low
+ 861.100000n V_low
+ 861.100001n V_low
+ 861.200000n V_low
+ 861.200001n V_low
+ 861.300000n V_low
+ 861.300001n V_low
+ 861.400000n V_low
+ 861.400001n V_low
+ 861.500000n V_low
+ 861.500001n V_low
+ 861.600000n V_low
+ 861.600001n V_low
+ 861.700000n V_low
+ 861.700001n V_low
+ 861.800000n V_low
+ 861.800001n V_low
+ 861.900000n V_low
+ 861.900001n V_low
+ 862.000000n V_low
+ 862.000001n V_hig
+ 862.100000n V_hig
+ 862.100001n V_hig
+ 862.200000n V_hig
+ 862.200001n V_hig
+ 862.300000n V_hig
+ 862.300001n V_hig
+ 862.400000n V_hig
+ 862.400001n V_hig
+ 862.500000n V_hig
+ 862.500001n V_hig
+ 862.600000n V_hig
+ 862.600001n V_hig
+ 862.700000n V_hig
+ 862.700001n V_hig
+ 862.800000n V_hig
+ 862.800001n V_hig
+ 862.900000n V_hig
+ 862.900001n V_hig
+ 863.000000n V_hig
+ 863.000001n V_low
+ 863.100000n V_low
+ 863.100001n V_low
+ 863.200000n V_low
+ 863.200001n V_low
+ 863.300000n V_low
+ 863.300001n V_low
+ 863.400000n V_low
+ 863.400001n V_low
+ 863.500000n V_low
+ 863.500001n V_low
+ 863.600000n V_low
+ 863.600001n V_low
+ 863.700000n V_low
+ 863.700001n V_low
+ 863.800000n V_low
+ 863.800001n V_low
+ 863.900000n V_low
+ 863.900001n V_low
+ 864.000000n V_low
+ 864.000001n V_hig
+ 864.100000n V_hig
+ 864.100001n V_hig
+ 864.200000n V_hig
+ 864.200001n V_hig
+ 864.300000n V_hig
+ 864.300001n V_hig
+ 864.400000n V_hig
+ 864.400001n V_hig
+ 864.500000n V_hig
+ 864.500001n V_hig
+ 864.600000n V_hig
+ 864.600001n V_hig
+ 864.700000n V_hig
+ 864.700001n V_hig
+ 864.800000n V_hig
+ 864.800001n V_hig
+ 864.900000n V_hig
+ 864.900001n V_hig
+ 865.000000n V_hig
+ 865.000001n V_hig
+ 865.100000n V_hig
+ 865.100001n V_hig
+ 865.200000n V_hig
+ 865.200001n V_hig
+ 865.300000n V_hig
+ 865.300001n V_hig
+ 865.400000n V_hig
+ 865.400001n V_hig
+ 865.500000n V_hig
+ 865.500001n V_hig
+ 865.600000n V_hig
+ 865.600001n V_hig
+ 865.700000n V_hig
+ 865.700001n V_hig
+ 865.800000n V_hig
+ 865.800001n V_hig
+ 865.900000n V_hig
+ 865.900001n V_hig
+ 866.000000n V_hig
+ 866.000001n V_hig
+ 866.100000n V_hig
+ 866.100001n V_hig
+ 866.200000n V_hig
+ 866.200001n V_hig
+ 866.300000n V_hig
+ 866.300001n V_hig
+ 866.400000n V_hig
+ 866.400001n V_hig
+ 866.500000n V_hig
+ 866.500001n V_hig
+ 866.600000n V_hig
+ 866.600001n V_hig
+ 866.700000n V_hig
+ 866.700001n V_hig
+ 866.800000n V_hig
+ 866.800001n V_hig
+ 866.900000n V_hig
+ 866.900001n V_hig
+ 867.000000n V_hig
+ 867.000001n V_low
+ 867.100000n V_low
+ 867.100001n V_low
+ 867.200000n V_low
+ 867.200001n V_low
+ 867.300000n V_low
+ 867.300001n V_low
+ 867.400000n V_low
+ 867.400001n V_low
+ 867.500000n V_low
+ 867.500001n V_low
+ 867.600000n V_low
+ 867.600001n V_low
+ 867.700000n V_low
+ 867.700001n V_low
+ 867.800000n V_low
+ 867.800001n V_low
+ 867.900000n V_low
+ 867.900001n V_low
+ 868.000000n V_low
+ 868.000001n V_low
+ 868.100000n V_low
+ 868.100001n V_low
+ 868.200000n V_low
+ 868.200001n V_low
+ 868.300000n V_low
+ 868.300001n V_low
+ 868.400000n V_low
+ 868.400001n V_low
+ 868.500000n V_low
+ 868.500001n V_low
+ 868.600000n V_low
+ 868.600001n V_low
+ 868.700000n V_low
+ 868.700001n V_low
+ 868.800000n V_low
+ 868.800001n V_low
+ 868.900000n V_low
+ 868.900001n V_low
+ 869.000000n V_low
+ 869.000001n V_hig
+ 869.100000n V_hig
+ 869.100001n V_hig
+ 869.200000n V_hig
+ 869.200001n V_hig
+ 869.300000n V_hig
+ 869.300001n V_hig
+ 869.400000n V_hig
+ 869.400001n V_hig
+ 869.500000n V_hig
+ 869.500001n V_hig
+ 869.600000n V_hig
+ 869.600001n V_hig
+ 869.700000n V_hig
+ 869.700001n V_hig
+ 869.800000n V_hig
+ 869.800001n V_hig
+ 869.900000n V_hig
+ 869.900001n V_hig
+ 870.000000n V_hig
+ 870.000001n V_low
+ 870.100000n V_low
+ 870.100001n V_low
+ 870.200000n V_low
+ 870.200001n V_low
+ 870.300000n V_low
+ 870.300001n V_low
+ 870.400000n V_low
+ 870.400001n V_low
+ 870.500000n V_low
+ 870.500001n V_low
+ 870.600000n V_low
+ 870.600001n V_low
+ 870.700000n V_low
+ 870.700001n V_low
+ 870.800000n V_low
+ 870.800001n V_low
+ 870.900000n V_low
+ 870.900001n V_low
+ 871.000000n V_low
+ 871.000001n V_hig
+ 871.100000n V_hig
+ 871.100001n V_hig
+ 871.200000n V_hig
+ 871.200001n V_hig
+ 871.300000n V_hig
+ 871.300001n V_hig
+ 871.400000n V_hig
+ 871.400001n V_hig
+ 871.500000n V_hig
+ 871.500001n V_hig
+ 871.600000n V_hig
+ 871.600001n V_hig
+ 871.700000n V_hig
+ 871.700001n V_hig
+ 871.800000n V_hig
+ 871.800001n V_hig
+ 871.900000n V_hig
+ 871.900001n V_hig
+ 872.000000n V_hig
+ 872.000001n V_low
+ 872.100000n V_low
+ 872.100001n V_low
+ 872.200000n V_low
+ 872.200001n V_low
+ 872.300000n V_low
+ 872.300001n V_low
+ 872.400000n V_low
+ 872.400001n V_low
+ 872.500000n V_low
+ 872.500001n V_low
+ 872.600000n V_low
+ 872.600001n V_low
+ 872.700000n V_low
+ 872.700001n V_low
+ 872.800000n V_low
+ 872.800001n V_low
+ 872.900000n V_low
+ 872.900001n V_low
+ 873.000000n V_low
+ 873.000001n V_low
+ 873.100000n V_low
+ 873.100001n V_low
+ 873.200000n V_low
+ 873.200001n V_low
+ 873.300000n V_low
+ 873.300001n V_low
+ 873.400000n V_low
+ 873.400001n V_low
+ 873.500000n V_low
+ 873.500001n V_low
+ 873.600000n V_low
+ 873.600001n V_low
+ 873.700000n V_low
+ 873.700001n V_low
+ 873.800000n V_low
+ 873.800001n V_low
+ 873.900000n V_low
+ 873.900001n V_low
+ 874.000000n V_low
+ 874.000001n V_hig
+ 874.100000n V_hig
+ 874.100001n V_hig
+ 874.200000n V_hig
+ 874.200001n V_hig
+ 874.300000n V_hig
+ 874.300001n V_hig
+ 874.400000n V_hig
+ 874.400001n V_hig
+ 874.500000n V_hig
+ 874.500001n V_hig
+ 874.600000n V_hig
+ 874.600001n V_hig
+ 874.700000n V_hig
+ 874.700001n V_hig
+ 874.800000n V_hig
+ 874.800001n V_hig
+ 874.900000n V_hig
+ 874.900001n V_hig
+ 875.000000n V_hig
+ 875.000001n V_hig
+ 875.100000n V_hig
+ 875.100001n V_hig
+ 875.200000n V_hig
+ 875.200001n V_hig
+ 875.300000n V_hig
+ 875.300001n V_hig
+ 875.400000n V_hig
+ 875.400001n V_hig
+ 875.500000n V_hig
+ 875.500001n V_hig
+ 875.600000n V_hig
+ 875.600001n V_hig
+ 875.700000n V_hig
+ 875.700001n V_hig
+ 875.800000n V_hig
+ 875.800001n V_hig
+ 875.900000n V_hig
+ 875.900001n V_hig
+ 876.000000n V_hig
+ 876.000001n V_hig
+ 876.100000n V_hig
+ 876.100001n V_hig
+ 876.200000n V_hig
+ 876.200001n V_hig
+ 876.300000n V_hig
+ 876.300001n V_hig
+ 876.400000n V_hig
+ 876.400001n V_hig
+ 876.500000n V_hig
+ 876.500001n V_hig
+ 876.600000n V_hig
+ 876.600001n V_hig
+ 876.700000n V_hig
+ 876.700001n V_hig
+ 876.800000n V_hig
+ 876.800001n V_hig
+ 876.900000n V_hig
+ 876.900001n V_hig
+ 877.000000n V_hig
+ 877.000001n V_low
+ 877.100000n V_low
+ 877.100001n V_low
+ 877.200000n V_low
+ 877.200001n V_low
+ 877.300000n V_low
+ 877.300001n V_low
+ 877.400000n V_low
+ 877.400001n V_low
+ 877.500000n V_low
+ 877.500001n V_low
+ 877.600000n V_low
+ 877.600001n V_low
+ 877.700000n V_low
+ 877.700001n V_low
+ 877.800000n V_low
+ 877.800001n V_low
+ 877.900000n V_low
+ 877.900001n V_low
+ 878.000000n V_low
+ 878.000001n V_low
+ 878.100000n V_low
+ 878.100001n V_low
+ 878.200000n V_low
+ 878.200001n V_low
+ 878.300000n V_low
+ 878.300001n V_low
+ 878.400000n V_low
+ 878.400001n V_low
+ 878.500000n V_low
+ 878.500001n V_low
+ 878.600000n V_low
+ 878.600001n V_low
+ 878.700000n V_low
+ 878.700001n V_low
+ 878.800000n V_low
+ 878.800001n V_low
+ 878.900000n V_low
+ 878.900001n V_low
+ 879.000000n V_low
+ 879.000001n V_hig
+ 879.100000n V_hig
+ 879.100001n V_hig
+ 879.200000n V_hig
+ 879.200001n V_hig
+ 879.300000n V_hig
+ 879.300001n V_hig
+ 879.400000n V_hig
+ 879.400001n V_hig
+ 879.500000n V_hig
+ 879.500001n V_hig
+ 879.600000n V_hig
+ 879.600001n V_hig
+ 879.700000n V_hig
+ 879.700001n V_hig
+ 879.800000n V_hig
+ 879.800001n V_hig
+ 879.900000n V_hig
+ 879.900001n V_hig
+ 880.000000n V_hig
+ 880.000001n V_low
+ 880.100000n V_low
+ 880.100001n V_low
+ 880.200000n V_low
+ 880.200001n V_low
+ 880.300000n V_low
+ 880.300001n V_low
+ 880.400000n V_low
+ 880.400001n V_low
+ 880.500000n V_low
+ 880.500001n V_low
+ 880.600000n V_low
+ 880.600001n V_low
+ 880.700000n V_low
+ 880.700001n V_low
+ 880.800000n V_low
+ 880.800001n V_low
+ 880.900000n V_low
+ 880.900001n V_low
+ 881.000000n V_low
+ 881.000001n V_low
+ 881.100000n V_low
+ 881.100001n V_low
+ 881.200000n V_low
+ 881.200001n V_low
+ 881.300000n V_low
+ 881.300001n V_low
+ 881.400000n V_low
+ 881.400001n V_low
+ 881.500000n V_low
+ 881.500001n V_low
+ 881.600000n V_low
+ 881.600001n V_low
+ 881.700000n V_low
+ 881.700001n V_low
+ 881.800000n V_low
+ 881.800001n V_low
+ 881.900000n V_low
+ 881.900001n V_low
+ 882.000000n V_low
+ 882.000001n V_hig
+ 882.100000n V_hig
+ 882.100001n V_hig
+ 882.200000n V_hig
+ 882.200001n V_hig
+ 882.300000n V_hig
+ 882.300001n V_hig
+ 882.400000n V_hig
+ 882.400001n V_hig
+ 882.500000n V_hig
+ 882.500001n V_hig
+ 882.600000n V_hig
+ 882.600001n V_hig
+ 882.700000n V_hig
+ 882.700001n V_hig
+ 882.800000n V_hig
+ 882.800001n V_hig
+ 882.900000n V_hig
+ 882.900001n V_hig
+ 883.000000n V_hig
+ 883.000001n V_hig
+ 883.100000n V_hig
+ 883.100001n V_hig
+ 883.200000n V_hig
+ 883.200001n V_hig
+ 883.300000n V_hig
+ 883.300001n V_hig
+ 883.400000n V_hig
+ 883.400001n V_hig
+ 883.500000n V_hig
+ 883.500001n V_hig
+ 883.600000n V_hig
+ 883.600001n V_hig
+ 883.700000n V_hig
+ 883.700001n V_hig
+ 883.800000n V_hig
+ 883.800001n V_hig
+ 883.900000n V_hig
+ 883.900001n V_hig
+ 884.000000n V_hig
+ 884.000001n V_hig
+ 884.100000n V_hig
+ 884.100001n V_hig
+ 884.200000n V_hig
+ 884.200001n V_hig
+ 884.300000n V_hig
+ 884.300001n V_hig
+ 884.400000n V_hig
+ 884.400001n V_hig
+ 884.500000n V_hig
+ 884.500001n V_hig
+ 884.600000n V_hig
+ 884.600001n V_hig
+ 884.700000n V_hig
+ 884.700001n V_hig
+ 884.800000n V_hig
+ 884.800001n V_hig
+ 884.900000n V_hig
+ 884.900001n V_hig
+ 885.000000n V_hig
+ 885.000001n V_hig
+ 885.100000n V_hig
+ 885.100001n V_hig
+ 885.200000n V_hig
+ 885.200001n V_hig
+ 885.300000n V_hig
+ 885.300001n V_hig
+ 885.400000n V_hig
+ 885.400001n V_hig
+ 885.500000n V_hig
+ 885.500001n V_hig
+ 885.600000n V_hig
+ 885.600001n V_hig
+ 885.700000n V_hig
+ 885.700001n V_hig
+ 885.800000n V_hig
+ 885.800001n V_hig
+ 885.900000n V_hig
+ 885.900001n V_hig
+ 886.000000n V_hig
+ 886.000001n V_low
+ 886.100000n V_low
+ 886.100001n V_low
+ 886.200000n V_low
+ 886.200001n V_low
+ 886.300000n V_low
+ 886.300001n V_low
+ 886.400000n V_low
+ 886.400001n V_low
+ 886.500000n V_low
+ 886.500001n V_low
+ 886.600000n V_low
+ 886.600001n V_low
+ 886.700000n V_low
+ 886.700001n V_low
+ 886.800000n V_low
+ 886.800001n V_low
+ 886.900000n V_low
+ 886.900001n V_low
+ 887.000000n V_low
+ 887.000001n V_hig
+ 887.100000n V_hig
+ 887.100001n V_hig
+ 887.200000n V_hig
+ 887.200001n V_hig
+ 887.300000n V_hig
+ 887.300001n V_hig
+ 887.400000n V_hig
+ 887.400001n V_hig
+ 887.500000n V_hig
+ 887.500001n V_hig
+ 887.600000n V_hig
+ 887.600001n V_hig
+ 887.700000n V_hig
+ 887.700001n V_hig
+ 887.800000n V_hig
+ 887.800001n V_hig
+ 887.900000n V_hig
+ 887.900001n V_hig
+ 888.000000n V_hig
+ 888.000001n V_hig
+ 888.100000n V_hig
+ 888.100001n V_hig
+ 888.200000n V_hig
+ 888.200001n V_hig
+ 888.300000n V_hig
+ 888.300001n V_hig
+ 888.400000n V_hig
+ 888.400001n V_hig
+ 888.500000n V_hig
+ 888.500001n V_hig
+ 888.600000n V_hig
+ 888.600001n V_hig
+ 888.700000n V_hig
+ 888.700001n V_hig
+ 888.800000n V_hig
+ 888.800001n V_hig
+ 888.900000n V_hig
+ 888.900001n V_hig
+ 889.000000n V_hig
+ 889.000001n V_low
+ 889.100000n V_low
+ 889.100001n V_low
+ 889.200000n V_low
+ 889.200001n V_low
+ 889.300000n V_low
+ 889.300001n V_low
+ 889.400000n V_low
+ 889.400001n V_low
+ 889.500000n V_low
+ 889.500001n V_low
+ 889.600000n V_low
+ 889.600001n V_low
+ 889.700000n V_low
+ 889.700001n V_low
+ 889.800000n V_low
+ 889.800001n V_low
+ 889.900000n V_low
+ 889.900001n V_low
+ 890.000000n V_low
+ 890.000001n V_hig
+ 890.100000n V_hig
+ 890.100001n V_hig
+ 890.200000n V_hig
+ 890.200001n V_hig
+ 890.300000n V_hig
+ 890.300001n V_hig
+ 890.400000n V_hig
+ 890.400001n V_hig
+ 890.500000n V_hig
+ 890.500001n V_hig
+ 890.600000n V_hig
+ 890.600001n V_hig
+ 890.700000n V_hig
+ 890.700001n V_hig
+ 890.800000n V_hig
+ 890.800001n V_hig
+ 890.900000n V_hig
+ 890.900001n V_hig
+ 891.000000n V_hig
+ 891.000001n V_hig
+ 891.100000n V_hig
+ 891.100001n V_hig
+ 891.200000n V_hig
+ 891.200001n V_hig
+ 891.300000n V_hig
+ 891.300001n V_hig
+ 891.400000n V_hig
+ 891.400001n V_hig
+ 891.500000n V_hig
+ 891.500001n V_hig
+ 891.600000n V_hig
+ 891.600001n V_hig
+ 891.700000n V_hig
+ 891.700001n V_hig
+ 891.800000n V_hig
+ 891.800001n V_hig
+ 891.900000n V_hig
+ 891.900001n V_hig
+ 892.000000n V_hig
+ 892.000001n V_low
+ 892.100000n V_low
+ 892.100001n V_low
+ 892.200000n V_low
+ 892.200001n V_low
+ 892.300000n V_low
+ 892.300001n V_low
+ 892.400000n V_low
+ 892.400001n V_low
+ 892.500000n V_low
+ 892.500001n V_low
+ 892.600000n V_low
+ 892.600001n V_low
+ 892.700000n V_low
+ 892.700001n V_low
+ 892.800000n V_low
+ 892.800001n V_low
+ 892.900000n V_low
+ 892.900001n V_low
+ 893.000000n V_low
+ 893.000001n V_low
+ 893.100000n V_low
+ 893.100001n V_low
+ 893.200000n V_low
+ 893.200001n V_low
+ 893.300000n V_low
+ 893.300001n V_low
+ 893.400000n V_low
+ 893.400001n V_low
+ 893.500000n V_low
+ 893.500001n V_low
+ 893.600000n V_low
+ 893.600001n V_low
+ 893.700000n V_low
+ 893.700001n V_low
+ 893.800000n V_low
+ 893.800001n V_low
+ 893.900000n V_low
+ 893.900001n V_low
+ 894.000000n V_low
+ 894.000001n V_hig
+ 894.100000n V_hig
+ 894.100001n V_hig
+ 894.200000n V_hig
+ 894.200001n V_hig
+ 894.300000n V_hig
+ 894.300001n V_hig
+ 894.400000n V_hig
+ 894.400001n V_hig
+ 894.500000n V_hig
+ 894.500001n V_hig
+ 894.600000n V_hig
+ 894.600001n V_hig
+ 894.700000n V_hig
+ 894.700001n V_hig
+ 894.800000n V_hig
+ 894.800001n V_hig
+ 894.900000n V_hig
+ 894.900001n V_hig
+ 895.000000n V_hig
+ 895.000001n V_hig
+ 895.100000n V_hig
+ 895.100001n V_hig
+ 895.200000n V_hig
+ 895.200001n V_hig
+ 895.300000n V_hig
+ 895.300001n V_hig
+ 895.400000n V_hig
+ 895.400001n V_hig
+ 895.500000n V_hig
+ 895.500001n V_hig
+ 895.600000n V_hig
+ 895.600001n V_hig
+ 895.700000n V_hig
+ 895.700001n V_hig
+ 895.800000n V_hig
+ 895.800001n V_hig
+ 895.900000n V_hig
+ 895.900001n V_hig
+ 896.000000n V_hig
+ 896.000001n V_low
+ 896.100000n V_low
+ 896.100001n V_low
+ 896.200000n V_low
+ 896.200001n V_low
+ 896.300000n V_low
+ 896.300001n V_low
+ 896.400000n V_low
+ 896.400001n V_low
+ 896.500000n V_low
+ 896.500001n V_low
+ 896.600000n V_low
+ 896.600001n V_low
+ 896.700000n V_low
+ 896.700001n V_low
+ 896.800000n V_low
+ 896.800001n V_low
+ 896.900000n V_low
+ 896.900001n V_low
+ 897.000000n V_low
+ 897.000001n V_low
+ 897.100000n V_low
+ 897.100001n V_low
+ 897.200000n V_low
+ 897.200001n V_low
+ 897.300000n V_low
+ 897.300001n V_low
+ 897.400000n V_low
+ 897.400001n V_low
+ 897.500000n V_low
+ 897.500001n V_low
+ 897.600000n V_low
+ 897.600001n V_low
+ 897.700000n V_low
+ 897.700001n V_low
+ 897.800000n V_low
+ 897.800001n V_low
+ 897.900000n V_low
+ 897.900001n V_low
+ 898.000000n V_low
+ 898.000001n V_low
+ 898.100000n V_low
+ 898.100001n V_low
+ 898.200000n V_low
+ 898.200001n V_low
+ 898.300000n V_low
+ 898.300001n V_low
+ 898.400000n V_low
+ 898.400001n V_low
+ 898.500000n V_low
+ 898.500001n V_low
+ 898.600000n V_low
+ 898.600001n V_low
+ 898.700000n V_low
+ 898.700001n V_low
+ 898.800000n V_low
+ 898.800001n V_low
+ 898.900000n V_low
+ 898.900001n V_low
+ 899.000000n V_low
+ 899.000001n V_hig
+ 899.100000n V_hig
+ 899.100001n V_hig
+ 899.200000n V_hig
+ 899.200001n V_hig
+ 899.300000n V_hig
+ 899.300001n V_hig
+ 899.400000n V_hig
+ 899.400001n V_hig
+ 899.500000n V_hig
+ 899.500001n V_hig
+ 899.600000n V_hig
+ 899.600001n V_hig
+ 899.700000n V_hig
+ 899.700001n V_hig
+ 899.800000n V_hig
+ 899.800001n V_hig
+ 899.900000n V_hig
+ 899.900001n V_hig
+ 900.000000n V_hig
+ 900.000001n V_low
+ 900.100000n V_low
+ 900.100001n V_low
+ 900.200000n V_low
+ 900.200001n V_low
+ 900.300000n V_low
+ 900.300001n V_low
+ 900.400000n V_low
+ 900.400001n V_low
+ 900.500000n V_low
+ 900.500001n V_low
+ 900.600000n V_low
+ 900.600001n V_low
+ 900.700000n V_low
+ 900.700001n V_low
+ 900.800000n V_low
+ 900.800001n V_low
+ 900.900000n V_low
+ 900.900001n V_low
+ 901.000000n V_low
+ 901.000001n V_low
+ 901.100000n V_low
+ 901.100001n V_low
+ 901.200000n V_low
+ 901.200001n V_low
+ 901.300000n V_low
+ 901.300001n V_low
+ 901.400000n V_low
+ 901.400001n V_low
+ 901.500000n V_low
+ 901.500001n V_low
+ 901.600000n V_low
+ 901.600001n V_low
+ 901.700000n V_low
+ 901.700001n V_low
+ 901.800000n V_low
+ 901.800001n V_low
+ 901.900000n V_low
+ 901.900001n V_low
+ 902.000000n V_low
+ 902.000001n V_hig
+ 902.100000n V_hig
+ 902.100001n V_hig
+ 902.200000n V_hig
+ 902.200001n V_hig
+ 902.300000n V_hig
+ 902.300001n V_hig
+ 902.400000n V_hig
+ 902.400001n V_hig
+ 902.500000n V_hig
+ 902.500001n V_hig
+ 902.600000n V_hig
+ 902.600001n V_hig
+ 902.700000n V_hig
+ 902.700001n V_hig
+ 902.800000n V_hig
+ 902.800001n V_hig
+ 902.900000n V_hig
+ 902.900001n V_hig
+ 903.000000n V_hig
+ 903.000001n V_hig
+ 903.100000n V_hig
+ 903.100001n V_hig
+ 903.200000n V_hig
+ 903.200001n V_hig
+ 903.300000n V_hig
+ 903.300001n V_hig
+ 903.400000n V_hig
+ 903.400001n V_hig
+ 903.500000n V_hig
+ 903.500001n V_hig
+ 903.600000n V_hig
+ 903.600001n V_hig
+ 903.700000n V_hig
+ 903.700001n V_hig
+ 903.800000n V_hig
+ 903.800001n V_hig
+ 903.900000n V_hig
+ 903.900001n V_hig
+ 904.000000n V_hig
+ 904.000001n V_hig
+ 904.100000n V_hig
+ 904.100001n V_hig
+ 904.200000n V_hig
+ 904.200001n V_hig
+ 904.300000n V_hig
+ 904.300001n V_hig
+ 904.400000n V_hig
+ 904.400001n V_hig
+ 904.500000n V_hig
+ 904.500001n V_hig
+ 904.600000n V_hig
+ 904.600001n V_hig
+ 904.700000n V_hig
+ 904.700001n V_hig
+ 904.800000n V_hig
+ 904.800001n V_hig
+ 904.900000n V_hig
+ 904.900001n V_hig
+ 905.000000n V_hig
+ 905.000001n V_hig
+ 905.100000n V_hig
+ 905.100001n V_hig
+ 905.200000n V_hig
+ 905.200001n V_hig
+ 905.300000n V_hig
+ 905.300001n V_hig
+ 905.400000n V_hig
+ 905.400001n V_hig
+ 905.500000n V_hig
+ 905.500001n V_hig
+ 905.600000n V_hig
+ 905.600001n V_hig
+ 905.700000n V_hig
+ 905.700001n V_hig
+ 905.800000n V_hig
+ 905.800001n V_hig
+ 905.900000n V_hig
+ 905.900001n V_hig
+ 906.000000n V_hig
+ 906.000001n V_low
+ 906.100000n V_low
+ 906.100001n V_low
+ 906.200000n V_low
+ 906.200001n V_low
+ 906.300000n V_low
+ 906.300001n V_low
+ 906.400000n V_low
+ 906.400001n V_low
+ 906.500000n V_low
+ 906.500001n V_low
+ 906.600000n V_low
+ 906.600001n V_low
+ 906.700000n V_low
+ 906.700001n V_low
+ 906.800000n V_low
+ 906.800001n V_low
+ 906.900000n V_low
+ 906.900001n V_low
+ 907.000000n V_low
+ 907.000001n V_hig
+ 907.100000n V_hig
+ 907.100001n V_hig
+ 907.200000n V_hig
+ 907.200001n V_hig
+ 907.300000n V_hig
+ 907.300001n V_hig
+ 907.400000n V_hig
+ 907.400001n V_hig
+ 907.500000n V_hig
+ 907.500001n V_hig
+ 907.600000n V_hig
+ 907.600001n V_hig
+ 907.700000n V_hig
+ 907.700001n V_hig
+ 907.800000n V_hig
+ 907.800001n V_hig
+ 907.900000n V_hig
+ 907.900001n V_hig
+ 908.000000n V_hig
+ 908.000001n V_low
+ 908.100000n V_low
+ 908.100001n V_low
+ 908.200000n V_low
+ 908.200001n V_low
+ 908.300000n V_low
+ 908.300001n V_low
+ 908.400000n V_low
+ 908.400001n V_low
+ 908.500000n V_low
+ 908.500001n V_low
+ 908.600000n V_low
+ 908.600001n V_low
+ 908.700000n V_low
+ 908.700001n V_low
+ 908.800000n V_low
+ 908.800001n V_low
+ 908.900000n V_low
+ 908.900001n V_low
+ 909.000000n V_low
+ 909.000001n V_low
+ 909.100000n V_low
+ 909.100001n V_low
+ 909.200000n V_low
+ 909.200001n V_low
+ 909.300000n V_low
+ 909.300001n V_low
+ 909.400000n V_low
+ 909.400001n V_low
+ 909.500000n V_low
+ 909.500001n V_low
+ 909.600000n V_low
+ 909.600001n V_low
+ 909.700000n V_low
+ 909.700001n V_low
+ 909.800000n V_low
+ 909.800001n V_low
+ 909.900000n V_low
+ 909.900001n V_low
+ 910.000000n V_low
+ 910.000001n V_hig
+ 910.100000n V_hig
+ 910.100001n V_hig
+ 910.200000n V_hig
+ 910.200001n V_hig
+ 910.300000n V_hig
+ 910.300001n V_hig
+ 910.400000n V_hig
+ 910.400001n V_hig
+ 910.500000n V_hig
+ 910.500001n V_hig
+ 910.600000n V_hig
+ 910.600001n V_hig
+ 910.700000n V_hig
+ 910.700001n V_hig
+ 910.800000n V_hig
+ 910.800001n V_hig
+ 910.900000n V_hig
+ 910.900001n V_hig
+ 911.000000n V_hig
+ 911.000001n V_hig
+ 911.100000n V_hig
+ 911.100001n V_hig
+ 911.200000n V_hig
+ 911.200001n V_hig
+ 911.300000n V_hig
+ 911.300001n V_hig
+ 911.400000n V_hig
+ 911.400001n V_hig
+ 911.500000n V_hig
+ 911.500001n V_hig
+ 911.600000n V_hig
+ 911.600001n V_hig
+ 911.700000n V_hig
+ 911.700001n V_hig
+ 911.800000n V_hig
+ 911.800001n V_hig
+ 911.900000n V_hig
+ 911.900001n V_hig
+ 912.000000n V_hig
+ 912.000001n V_low
+ 912.100000n V_low
+ 912.100001n V_low
+ 912.200000n V_low
+ 912.200001n V_low
+ 912.300000n V_low
+ 912.300001n V_low
+ 912.400000n V_low
+ 912.400001n V_low
+ 912.500000n V_low
+ 912.500001n V_low
+ 912.600000n V_low
+ 912.600001n V_low
+ 912.700000n V_low
+ 912.700001n V_low
+ 912.800000n V_low
+ 912.800001n V_low
+ 912.900000n V_low
+ 912.900001n V_low
+ 913.000000n V_low
+ 913.000001n V_low
+ 913.100000n V_low
+ 913.100001n V_low
+ 913.200000n V_low
+ 913.200001n V_low
+ 913.300000n V_low
+ 913.300001n V_low
+ 913.400000n V_low
+ 913.400001n V_low
+ 913.500000n V_low
+ 913.500001n V_low
+ 913.600000n V_low
+ 913.600001n V_low
+ 913.700000n V_low
+ 913.700001n V_low
+ 913.800000n V_low
+ 913.800001n V_low
+ 913.900000n V_low
+ 913.900001n V_low
+ 914.000000n V_low
+ 914.000001n V_hig
+ 914.100000n V_hig
+ 914.100001n V_hig
+ 914.200000n V_hig
+ 914.200001n V_hig
+ 914.300000n V_hig
+ 914.300001n V_hig
+ 914.400000n V_hig
+ 914.400001n V_hig
+ 914.500000n V_hig
+ 914.500001n V_hig
+ 914.600000n V_hig
+ 914.600001n V_hig
+ 914.700000n V_hig
+ 914.700001n V_hig
+ 914.800000n V_hig
+ 914.800001n V_hig
+ 914.900000n V_hig
+ 914.900001n V_hig
+ 915.000000n V_hig
+ 915.000001n V_hig
+ 915.100000n V_hig
+ 915.100001n V_hig
+ 915.200000n V_hig
+ 915.200001n V_hig
+ 915.300000n V_hig
+ 915.300001n V_hig
+ 915.400000n V_hig
+ 915.400001n V_hig
+ 915.500000n V_hig
+ 915.500001n V_hig
+ 915.600000n V_hig
+ 915.600001n V_hig
+ 915.700000n V_hig
+ 915.700001n V_hig
+ 915.800000n V_hig
+ 915.800001n V_hig
+ 915.900000n V_hig
+ 915.900001n V_hig
+ 916.000000n V_hig
+ 916.000001n V_hig
+ 916.100000n V_hig
+ 916.100001n V_hig
+ 916.200000n V_hig
+ 916.200001n V_hig
+ 916.300000n V_hig
+ 916.300001n V_hig
+ 916.400000n V_hig
+ 916.400001n V_hig
+ 916.500000n V_hig
+ 916.500001n V_hig
+ 916.600000n V_hig
+ 916.600001n V_hig
+ 916.700000n V_hig
+ 916.700001n V_hig
+ 916.800000n V_hig
+ 916.800001n V_hig
+ 916.900000n V_hig
+ 916.900001n V_hig
+ 917.000000n V_hig
+ 917.000001n V_low
+ 917.100000n V_low
+ 917.100001n V_low
+ 917.200000n V_low
+ 917.200001n V_low
+ 917.300000n V_low
+ 917.300001n V_low
+ 917.400000n V_low
+ 917.400001n V_low
+ 917.500000n V_low
+ 917.500001n V_low
+ 917.600000n V_low
+ 917.600001n V_low
+ 917.700000n V_low
+ 917.700001n V_low
+ 917.800000n V_low
+ 917.800001n V_low
+ 917.900000n V_low
+ 917.900001n V_low
+ 918.000000n V_low
+ 918.000001n V_low
+ 918.100000n V_low
+ 918.100001n V_low
+ 918.200000n V_low
+ 918.200001n V_low
+ 918.300000n V_low
+ 918.300001n V_low
+ 918.400000n V_low
+ 918.400001n V_low
+ 918.500000n V_low
+ 918.500001n V_low
+ 918.600000n V_low
+ 918.600001n V_low
+ 918.700000n V_low
+ 918.700001n V_low
+ 918.800000n V_low
+ 918.800001n V_low
+ 918.900000n V_low
+ 918.900001n V_low
+ 919.000000n V_low
+ 919.000001n V_hig
+ 919.100000n V_hig
+ 919.100001n V_hig
+ 919.200000n V_hig
+ 919.200001n V_hig
+ 919.300000n V_hig
+ 919.300001n V_hig
+ 919.400000n V_hig
+ 919.400001n V_hig
+ 919.500000n V_hig
+ 919.500001n V_hig
+ 919.600000n V_hig
+ 919.600001n V_hig
+ 919.700000n V_hig
+ 919.700001n V_hig
+ 919.800000n V_hig
+ 919.800001n V_hig
+ 919.900000n V_hig
+ 919.900001n V_hig
+ 920.000000n V_hig
+ 920.000001n V_low
+ 920.100000n V_low
+ 920.100001n V_low
+ 920.200000n V_low
+ 920.200001n V_low
+ 920.300000n V_low
+ 920.300001n V_low
+ 920.400000n V_low
+ 920.400001n V_low
+ 920.500000n V_low
+ 920.500001n V_low
+ 920.600000n V_low
+ 920.600001n V_low
+ 920.700000n V_low
+ 920.700001n V_low
+ 920.800000n V_low
+ 920.800001n V_low
+ 920.900000n V_low
+ 920.900001n V_low
+ 921.000000n V_low
+ 921.000001n V_low
+ 921.100000n V_low
+ 921.100001n V_low
+ 921.200000n V_low
+ 921.200001n V_low
+ 921.300000n V_low
+ 921.300001n V_low
+ 921.400000n V_low
+ 921.400001n V_low
+ 921.500000n V_low
+ 921.500001n V_low
+ 921.600000n V_low
+ 921.600001n V_low
+ 921.700000n V_low
+ 921.700001n V_low
+ 921.800000n V_low
+ 921.800001n V_low
+ 921.900000n V_low
+ 921.900001n V_low
+ 922.000000n V_low
+ 922.000001n V_low
+ 922.100000n V_low
+ 922.100001n V_low
+ 922.200000n V_low
+ 922.200001n V_low
+ 922.300000n V_low
+ 922.300001n V_low
+ 922.400000n V_low
+ 922.400001n V_low
+ 922.500000n V_low
+ 922.500001n V_low
+ 922.600000n V_low
+ 922.600001n V_low
+ 922.700000n V_low
+ 922.700001n V_low
+ 922.800000n V_low
+ 922.800001n V_low
+ 922.900000n V_low
+ 922.900001n V_low
+ 923.000000n V_low
+ 923.000001n V_hig
+ 923.100000n V_hig
+ 923.100001n V_hig
+ 923.200000n V_hig
+ 923.200001n V_hig
+ 923.300000n V_hig
+ 923.300001n V_hig
+ 923.400000n V_hig
+ 923.400001n V_hig
+ 923.500000n V_hig
+ 923.500001n V_hig
+ 923.600000n V_hig
+ 923.600001n V_hig
+ 923.700000n V_hig
+ 923.700001n V_hig
+ 923.800000n V_hig
+ 923.800001n V_hig
+ 923.900000n V_hig
+ 923.900001n V_hig
+ 924.000000n V_hig
+ 924.000001n V_low
+ 924.100000n V_low
+ 924.100001n V_low
+ 924.200000n V_low
+ 924.200001n V_low
+ 924.300000n V_low
+ 924.300001n V_low
+ 924.400000n V_low
+ 924.400001n V_low
+ 924.500000n V_low
+ 924.500001n V_low
+ 924.600000n V_low
+ 924.600001n V_low
+ 924.700000n V_low
+ 924.700001n V_low
+ 924.800000n V_low
+ 924.800001n V_low
+ 924.900000n V_low
+ 924.900001n V_low
+ 925.000000n V_low
+ 925.000001n V_low
+ 925.100000n V_low
+ 925.100001n V_low
+ 925.200000n V_low
+ 925.200001n V_low
+ 925.300000n V_low
+ 925.300001n V_low
+ 925.400000n V_low
+ 925.400001n V_low
+ 925.500000n V_low
+ 925.500001n V_low
+ 925.600000n V_low
+ 925.600001n V_low
+ 925.700000n V_low
+ 925.700001n V_low
+ 925.800000n V_low
+ 925.800001n V_low
+ 925.900000n V_low
+ 925.900001n V_low
+ 926.000000n V_low
+ 926.000001n V_low
+ 926.100000n V_low
+ 926.100001n V_low
+ 926.200000n V_low
+ 926.200001n V_low
+ 926.300000n V_low
+ 926.300001n V_low
+ 926.400000n V_low
+ 926.400001n V_low
+ 926.500000n V_low
+ 926.500001n V_low
+ 926.600000n V_low
+ 926.600001n V_low
+ 926.700000n V_low
+ 926.700001n V_low
+ 926.800000n V_low
+ 926.800001n V_low
+ 926.900000n V_low
+ 926.900001n V_low
+ 927.000000n V_low
+ 927.000001n V_low
+ 927.100000n V_low
+ 927.100001n V_low
+ 927.200000n V_low
+ 927.200001n V_low
+ 927.300000n V_low
+ 927.300001n V_low
+ 927.400000n V_low
+ 927.400001n V_low
+ 927.500000n V_low
+ 927.500001n V_low
+ 927.600000n V_low
+ 927.600001n V_low
+ 927.700000n V_low
+ 927.700001n V_low
+ 927.800000n V_low
+ 927.800001n V_low
+ 927.900000n V_low
+ 927.900001n V_low
+ 928.000000n V_low
+ 928.000001n V_low
+ 928.100000n V_low
+ 928.100001n V_low
+ 928.200000n V_low
+ 928.200001n V_low
+ 928.300000n V_low
+ 928.300001n V_low
+ 928.400000n V_low
+ 928.400001n V_low
+ 928.500000n V_low
+ 928.500001n V_low
+ 928.600000n V_low
+ 928.600001n V_low
+ 928.700000n V_low
+ 928.700001n V_low
+ 928.800000n V_low
+ 928.800001n V_low
+ 928.900000n V_low
+ 928.900001n V_low
+ 929.000000n V_low
+ 929.000001n V_hig
+ 929.100000n V_hig
+ 929.100001n V_hig
+ 929.200000n V_hig
+ 929.200001n V_hig
+ 929.300000n V_hig
+ 929.300001n V_hig
+ 929.400000n V_hig
+ 929.400001n V_hig
+ 929.500000n V_hig
+ 929.500001n V_hig
+ 929.600000n V_hig
+ 929.600001n V_hig
+ 929.700000n V_hig
+ 929.700001n V_hig
+ 929.800000n V_hig
+ 929.800001n V_hig
+ 929.900000n V_hig
+ 929.900001n V_hig
+ 930.000000n V_hig
+ 930.000001n V_hig
+ 930.100000n V_hig
+ 930.100001n V_hig
+ 930.200000n V_hig
+ 930.200001n V_hig
+ 930.300000n V_hig
+ 930.300001n V_hig
+ 930.400000n V_hig
+ 930.400001n V_hig
+ 930.500000n V_hig
+ 930.500001n V_hig
+ 930.600000n V_hig
+ 930.600001n V_hig
+ 930.700000n V_hig
+ 930.700001n V_hig
+ 930.800000n V_hig
+ 930.800001n V_hig
+ 930.900000n V_hig
+ 930.900001n V_hig
+ 931.000000n V_hig
+ 931.000001n V_hig
+ 931.100000n V_hig
+ 931.100001n V_hig
+ 931.200000n V_hig
+ 931.200001n V_hig
+ 931.300000n V_hig
+ 931.300001n V_hig
+ 931.400000n V_hig
+ 931.400001n V_hig
+ 931.500000n V_hig
+ 931.500001n V_hig
+ 931.600000n V_hig
+ 931.600001n V_hig
+ 931.700000n V_hig
+ 931.700001n V_hig
+ 931.800000n V_hig
+ 931.800001n V_hig
+ 931.900000n V_hig
+ 931.900001n V_hig
+ 932.000000n V_hig
+ 932.000001n V_low
+ 932.100000n V_low
+ 932.100001n V_low
+ 932.200000n V_low
+ 932.200001n V_low
+ 932.300000n V_low
+ 932.300001n V_low
+ 932.400000n V_low
+ 932.400001n V_low
+ 932.500000n V_low
+ 932.500001n V_low
+ 932.600000n V_low
+ 932.600001n V_low
+ 932.700000n V_low
+ 932.700001n V_low
+ 932.800000n V_low
+ 932.800001n V_low
+ 932.900000n V_low
+ 932.900001n V_low
+ 933.000000n V_low
+ 933.000001n V_hig
+ 933.100000n V_hig
+ 933.100001n V_hig
+ 933.200000n V_hig
+ 933.200001n V_hig
+ 933.300000n V_hig
+ 933.300001n V_hig
+ 933.400000n V_hig
+ 933.400001n V_hig
+ 933.500000n V_hig
+ 933.500001n V_hig
+ 933.600000n V_hig
+ 933.600001n V_hig
+ 933.700000n V_hig
+ 933.700001n V_hig
+ 933.800000n V_hig
+ 933.800001n V_hig
+ 933.900000n V_hig
+ 933.900001n V_hig
+ 934.000000n V_hig
+ 934.000001n V_hig
+ 934.100000n V_hig
+ 934.100001n V_hig
+ 934.200000n V_hig
+ 934.200001n V_hig
+ 934.300000n V_hig
+ 934.300001n V_hig
+ 934.400000n V_hig
+ 934.400001n V_hig
+ 934.500000n V_hig
+ 934.500001n V_hig
+ 934.600000n V_hig
+ 934.600001n V_hig
+ 934.700000n V_hig
+ 934.700001n V_hig
+ 934.800000n V_hig
+ 934.800001n V_hig
+ 934.900000n V_hig
+ 934.900001n V_hig
+ 935.000000n V_hig
+ 935.000001n V_low
+ 935.100000n V_low
+ 935.100001n V_low
+ 935.200000n V_low
+ 935.200001n V_low
+ 935.300000n V_low
+ 935.300001n V_low
+ 935.400000n V_low
+ 935.400001n V_low
+ 935.500000n V_low
+ 935.500001n V_low
+ 935.600000n V_low
+ 935.600001n V_low
+ 935.700000n V_low
+ 935.700001n V_low
+ 935.800000n V_low
+ 935.800001n V_low
+ 935.900000n V_low
+ 935.900001n V_low
+ 936.000000n V_low
+ 936.000001n V_low
+ 936.100000n V_low
+ 936.100001n V_low
+ 936.200000n V_low
+ 936.200001n V_low
+ 936.300000n V_low
+ 936.300001n V_low
+ 936.400000n V_low
+ 936.400001n V_low
+ 936.500000n V_low
+ 936.500001n V_low
+ 936.600000n V_low
+ 936.600001n V_low
+ 936.700000n V_low
+ 936.700001n V_low
+ 936.800000n V_low
+ 936.800001n V_low
+ 936.900000n V_low
+ 936.900001n V_low
+ 937.000000n V_low
+ 937.000001n V_hig
+ 937.100000n V_hig
+ 937.100001n V_hig
+ 937.200000n V_hig
+ 937.200001n V_hig
+ 937.300000n V_hig
+ 937.300001n V_hig
+ 937.400000n V_hig
+ 937.400001n V_hig
+ 937.500000n V_hig
+ 937.500001n V_hig
+ 937.600000n V_hig
+ 937.600001n V_hig
+ 937.700000n V_hig
+ 937.700001n V_hig
+ 937.800000n V_hig
+ 937.800001n V_hig
+ 937.900000n V_hig
+ 937.900001n V_hig
+ 938.000000n V_hig
+ 938.000001n V_hig
+ 938.100000n V_hig
+ 938.100001n V_hig
+ 938.200000n V_hig
+ 938.200001n V_hig
+ 938.300000n V_hig
+ 938.300001n V_hig
+ 938.400000n V_hig
+ 938.400001n V_hig
+ 938.500000n V_hig
+ 938.500001n V_hig
+ 938.600000n V_hig
+ 938.600001n V_hig
+ 938.700000n V_hig
+ 938.700001n V_hig
+ 938.800000n V_hig
+ 938.800001n V_hig
+ 938.900000n V_hig
+ 938.900001n V_hig
+ 939.000000n V_hig
+ 939.000001n V_low
+ 939.100000n V_low
+ 939.100001n V_low
+ 939.200000n V_low
+ 939.200001n V_low
+ 939.300000n V_low
+ 939.300001n V_low
+ 939.400000n V_low
+ 939.400001n V_low
+ 939.500000n V_low
+ 939.500001n V_low
+ 939.600000n V_low
+ 939.600001n V_low
+ 939.700000n V_low
+ 939.700001n V_low
+ 939.800000n V_low
+ 939.800001n V_low
+ 939.900000n V_low
+ 939.900001n V_low
+ 940.000000n V_low
+ 940.000001n V_hig
+ 940.100000n V_hig
+ 940.100001n V_hig
+ 940.200000n V_hig
+ 940.200001n V_hig
+ 940.300000n V_hig
+ 940.300001n V_hig
+ 940.400000n V_hig
+ 940.400001n V_hig
+ 940.500000n V_hig
+ 940.500001n V_hig
+ 940.600000n V_hig
+ 940.600001n V_hig
+ 940.700000n V_hig
+ 940.700001n V_hig
+ 940.800000n V_hig
+ 940.800001n V_hig
+ 940.900000n V_hig
+ 940.900001n V_hig
+ 941.000000n V_hig
+ 941.000001n V_hig
+ 941.100000n V_hig
+ 941.100001n V_hig
+ 941.200000n V_hig
+ 941.200001n V_hig
+ 941.300000n V_hig
+ 941.300001n V_hig
+ 941.400000n V_hig
+ 941.400001n V_hig
+ 941.500000n V_hig
+ 941.500001n V_hig
+ 941.600000n V_hig
+ 941.600001n V_hig
+ 941.700000n V_hig
+ 941.700001n V_hig
+ 941.800000n V_hig
+ 941.800001n V_hig
+ 941.900000n V_hig
+ 941.900001n V_hig
+ 942.000000n V_hig
+ 942.000001n V_hig
+ 942.100000n V_hig
+ 942.100001n V_hig
+ 942.200000n V_hig
+ 942.200001n V_hig
+ 942.300000n V_hig
+ 942.300001n V_hig
+ 942.400000n V_hig
+ 942.400001n V_hig
+ 942.500000n V_hig
+ 942.500001n V_hig
+ 942.600000n V_hig
+ 942.600001n V_hig
+ 942.700000n V_hig
+ 942.700001n V_hig
+ 942.800000n V_hig
+ 942.800001n V_hig
+ 942.900000n V_hig
+ 942.900001n V_hig
+ 943.000000n V_hig
+ 943.000001n V_hig
+ 943.100000n V_hig
+ 943.100001n V_hig
+ 943.200000n V_hig
+ 943.200001n V_hig
+ 943.300000n V_hig
+ 943.300001n V_hig
+ 943.400000n V_hig
+ 943.400001n V_hig
+ 943.500000n V_hig
+ 943.500001n V_hig
+ 943.600000n V_hig
+ 943.600001n V_hig
+ 943.700000n V_hig
+ 943.700001n V_hig
+ 943.800000n V_hig
+ 943.800001n V_hig
+ 943.900000n V_hig
+ 943.900001n V_hig
+ 944.000000n V_hig
+ 944.000001n V_low
+ 944.100000n V_low
+ 944.100001n V_low
+ 944.200000n V_low
+ 944.200001n V_low
+ 944.300000n V_low
+ 944.300001n V_low
+ 944.400000n V_low
+ 944.400001n V_low
+ 944.500000n V_low
+ 944.500001n V_low
+ 944.600000n V_low
+ 944.600001n V_low
+ 944.700000n V_low
+ 944.700001n V_low
+ 944.800000n V_low
+ 944.800001n V_low
+ 944.900000n V_low
+ 944.900001n V_low
+ 945.000000n V_low
+ 945.000001n V_hig
+ 945.100000n V_hig
+ 945.100001n V_hig
+ 945.200000n V_hig
+ 945.200001n V_hig
+ 945.300000n V_hig
+ 945.300001n V_hig
+ 945.400000n V_hig
+ 945.400001n V_hig
+ 945.500000n V_hig
+ 945.500001n V_hig
+ 945.600000n V_hig
+ 945.600001n V_hig
+ 945.700000n V_hig
+ 945.700001n V_hig
+ 945.800000n V_hig
+ 945.800001n V_hig
+ 945.900000n V_hig
+ 945.900001n V_hig
+ 946.000000n V_hig
+ 946.000001n V_hig
+ 946.100000n V_hig
+ 946.100001n V_hig
+ 946.200000n V_hig
+ 946.200001n V_hig
+ 946.300000n V_hig
+ 946.300001n V_hig
+ 946.400000n V_hig
+ 946.400001n V_hig
+ 946.500000n V_hig
+ 946.500001n V_hig
+ 946.600000n V_hig
+ 946.600001n V_hig
+ 946.700000n V_hig
+ 946.700001n V_hig
+ 946.800000n V_hig
+ 946.800001n V_hig
+ 946.900000n V_hig
+ 946.900001n V_hig
+ 947.000000n V_hig
+ 947.000001n V_hig
+ 947.100000n V_hig
+ 947.100001n V_hig
+ 947.200000n V_hig
+ 947.200001n V_hig
+ 947.300000n V_hig
+ 947.300001n V_hig
+ 947.400000n V_hig
+ 947.400001n V_hig
+ 947.500000n V_hig
+ 947.500001n V_hig
+ 947.600000n V_hig
+ 947.600001n V_hig
+ 947.700000n V_hig
+ 947.700001n V_hig
+ 947.800000n V_hig
+ 947.800001n V_hig
+ 947.900000n V_hig
+ 947.900001n V_hig
+ 948.000000n V_hig
+ 948.000001n V_low
+ 948.100000n V_low
+ 948.100001n V_low
+ 948.200000n V_low
+ 948.200001n V_low
+ 948.300000n V_low
+ 948.300001n V_low
+ 948.400000n V_low
+ 948.400001n V_low
+ 948.500000n V_low
+ 948.500001n V_low
+ 948.600000n V_low
+ 948.600001n V_low
+ 948.700000n V_low
+ 948.700001n V_low
+ 948.800000n V_low
+ 948.800001n V_low
+ 948.900000n V_low
+ 948.900001n V_low
+ 949.000000n V_low
+ 949.000001n V_hig
+ 949.100000n V_hig
+ 949.100001n V_hig
+ 949.200000n V_hig
+ 949.200001n V_hig
+ 949.300000n V_hig
+ 949.300001n V_hig
+ 949.400000n V_hig
+ 949.400001n V_hig
+ 949.500000n V_hig
+ 949.500001n V_hig
+ 949.600000n V_hig
+ 949.600001n V_hig
+ 949.700000n V_hig
+ 949.700001n V_hig
+ 949.800000n V_hig
+ 949.800001n V_hig
+ 949.900000n V_hig
+ 949.900001n V_hig
+ 950.000000n V_hig
+ 950.000001n V_hig
+ 950.100000n V_hig
+ 950.100001n V_hig
+ 950.200000n V_hig
+ 950.200001n V_hig
+ 950.300000n V_hig
+ 950.300001n V_hig
+ 950.400000n V_hig
+ 950.400001n V_hig
+ 950.500000n V_hig
+ 950.500001n V_hig
+ 950.600000n V_hig
+ 950.600001n V_hig
+ 950.700000n V_hig
+ 950.700001n V_hig
+ 950.800000n V_hig
+ 950.800001n V_hig
+ 950.900000n V_hig
+ 950.900001n V_hig
+ 951.000000n V_hig
+ 951.000001n V_hig
+ 951.100000n V_hig
+ 951.100001n V_hig
+ 951.200000n V_hig
+ 951.200001n V_hig
+ 951.300000n V_hig
+ 951.300001n V_hig
+ 951.400000n V_hig
+ 951.400001n V_hig
+ 951.500000n V_hig
+ 951.500001n V_hig
+ 951.600000n V_hig
+ 951.600001n V_hig
+ 951.700000n V_hig
+ 951.700001n V_hig
+ 951.800000n V_hig
+ 951.800001n V_hig
+ 951.900000n V_hig
+ 951.900001n V_hig
+ 952.000000n V_hig
+ 952.000001n V_hig
+ 952.100000n V_hig
+ 952.100001n V_hig
+ 952.200000n V_hig
+ 952.200001n V_hig
+ 952.300000n V_hig
+ 952.300001n V_hig
+ 952.400000n V_hig
+ 952.400001n V_hig
+ 952.500000n V_hig
+ 952.500001n V_hig
+ 952.600000n V_hig
+ 952.600001n V_hig
+ 952.700000n V_hig
+ 952.700001n V_hig
+ 952.800000n V_hig
+ 952.800001n V_hig
+ 952.900000n V_hig
+ 952.900001n V_hig
+ 953.000000n V_hig
+ 953.000001n V_hig
+ 953.100000n V_hig
+ 953.100001n V_hig
+ 953.200000n V_hig
+ 953.200001n V_hig
+ 953.300000n V_hig
+ 953.300001n V_hig
+ 953.400000n V_hig
+ 953.400001n V_hig
+ 953.500000n V_hig
+ 953.500001n V_hig
+ 953.600000n V_hig
+ 953.600001n V_hig
+ 953.700000n V_hig
+ 953.700001n V_hig
+ 953.800000n V_hig
+ 953.800001n V_hig
+ 953.900000n V_hig
+ 953.900001n V_hig
+ 954.000000n V_hig
+ 954.000001n V_hig
+ 954.100000n V_hig
+ 954.100001n V_hig
+ 954.200000n V_hig
+ 954.200001n V_hig
+ 954.300000n V_hig
+ 954.300001n V_hig
+ 954.400000n V_hig
+ 954.400001n V_hig
+ 954.500000n V_hig
+ 954.500001n V_hig
+ 954.600000n V_hig
+ 954.600001n V_hig
+ 954.700000n V_hig
+ 954.700001n V_hig
+ 954.800000n V_hig
+ 954.800001n V_hig
+ 954.900000n V_hig
+ 954.900001n V_hig
+ 955.000000n V_hig
+ 955.000001n V_hig
+ 955.100000n V_hig
+ 955.100001n V_hig
+ 955.200000n V_hig
+ 955.200001n V_hig
+ 955.300000n V_hig
+ 955.300001n V_hig
+ 955.400000n V_hig
+ 955.400001n V_hig
+ 955.500000n V_hig
+ 955.500001n V_hig
+ 955.600000n V_hig
+ 955.600001n V_hig
+ 955.700000n V_hig
+ 955.700001n V_hig
+ 955.800000n V_hig
+ 955.800001n V_hig
+ 955.900000n V_hig
+ 955.900001n V_hig
+ 956.000000n V_hig
+ 956.000001n V_hig
+ 956.100000n V_hig
+ 956.100001n V_hig
+ 956.200000n V_hig
+ 956.200001n V_hig
+ 956.300000n V_hig
+ 956.300001n V_hig
+ 956.400000n V_hig
+ 956.400001n V_hig
+ 956.500000n V_hig
+ 956.500001n V_hig
+ 956.600000n V_hig
+ 956.600001n V_hig
+ 956.700000n V_hig
+ 956.700001n V_hig
+ 956.800000n V_hig
+ 956.800001n V_hig
+ 956.900000n V_hig
+ 956.900001n V_hig
+ 957.000000n V_hig
+ 957.000001n V_hig
+ 957.100000n V_hig
+ 957.100001n V_hig
+ 957.200000n V_hig
+ 957.200001n V_hig
+ 957.300000n V_hig
+ 957.300001n V_hig
+ 957.400000n V_hig
+ 957.400001n V_hig
+ 957.500000n V_hig
+ 957.500001n V_hig
+ 957.600000n V_hig
+ 957.600001n V_hig
+ 957.700000n V_hig
+ 957.700001n V_hig
+ 957.800000n V_hig
+ 957.800001n V_hig
+ 957.900000n V_hig
+ 957.900001n V_hig
+ 958.000000n V_hig
+ 958.000001n V_low
+ 958.100000n V_low
+ 958.100001n V_low
+ 958.200000n V_low
+ 958.200001n V_low
+ 958.300000n V_low
+ 958.300001n V_low
+ 958.400000n V_low
+ 958.400001n V_low
+ 958.500000n V_low
+ 958.500001n V_low
+ 958.600000n V_low
+ 958.600001n V_low
+ 958.700000n V_low
+ 958.700001n V_low
+ 958.800000n V_low
+ 958.800001n V_low
+ 958.900000n V_low
+ 958.900001n V_low
+ 959.000000n V_low
+ 959.000001n V_low
+ 959.100000n V_low
+ 959.100001n V_low
+ 959.200000n V_low
+ 959.200001n V_low
+ 959.300000n V_low
+ 959.300001n V_low
+ 959.400000n V_low
+ 959.400001n V_low
+ 959.500000n V_low
+ 959.500001n V_low
+ 959.600000n V_low
+ 959.600001n V_low
+ 959.700000n V_low
+ 959.700001n V_low
+ 959.800000n V_low
+ 959.800001n V_low
+ 959.900000n V_low
+ 959.900001n V_low
+ 960.000000n V_low
+ 960.000001n V_low
+ 960.100000n V_low
+ 960.100001n V_low
+ 960.200000n V_low
+ 960.200001n V_low
+ 960.300000n V_low
+ 960.300001n V_low
+ 960.400000n V_low
+ 960.400001n V_low
+ 960.500000n V_low
+ 960.500001n V_low
+ 960.600000n V_low
+ 960.600001n V_low
+ 960.700000n V_low
+ 960.700001n V_low
+ 960.800000n V_low
+ 960.800001n V_low
+ 960.900000n V_low
+ 960.900001n V_low
+ 961.000000n V_low
+ 961.000001n V_hig
+ 961.100000n V_hig
+ 961.100001n V_hig
+ 961.200000n V_hig
+ 961.200001n V_hig
+ 961.300000n V_hig
+ 961.300001n V_hig
+ 961.400000n V_hig
+ 961.400001n V_hig
+ 961.500000n V_hig
+ 961.500001n V_hig
+ 961.600000n V_hig
+ 961.600001n V_hig
+ 961.700000n V_hig
+ 961.700001n V_hig
+ 961.800000n V_hig
+ 961.800001n V_hig
+ 961.900000n V_hig
+ 961.900001n V_hig
+ 962.000000n V_hig
+ 962.000001n V_low
+ 962.100000n V_low
+ 962.100001n V_low
+ 962.200000n V_low
+ 962.200001n V_low
+ 962.300000n V_low
+ 962.300001n V_low
+ 962.400000n V_low
+ 962.400001n V_low
+ 962.500000n V_low
+ 962.500001n V_low
+ 962.600000n V_low
+ 962.600001n V_low
+ 962.700000n V_low
+ 962.700001n V_low
+ 962.800000n V_low
+ 962.800001n V_low
+ 962.900000n V_low
+ 962.900001n V_low
+ 963.000000n V_low
+ 963.000001n V_hig
+ 963.100000n V_hig
+ 963.100001n V_hig
+ 963.200000n V_hig
+ 963.200001n V_hig
+ 963.300000n V_hig
+ 963.300001n V_hig
+ 963.400000n V_hig
+ 963.400001n V_hig
+ 963.500000n V_hig
+ 963.500001n V_hig
+ 963.600000n V_hig
+ 963.600001n V_hig
+ 963.700000n V_hig
+ 963.700001n V_hig
+ 963.800000n V_hig
+ 963.800001n V_hig
+ 963.900000n V_hig
+ 963.900001n V_hig
+ 964.000000n V_hig
+ 964.000001n V_hig
+ 964.100000n V_hig
+ 964.100001n V_hig
+ 964.200000n V_hig
+ 964.200001n V_hig
+ 964.300000n V_hig
+ 964.300001n V_hig
+ 964.400000n V_hig
+ 964.400001n V_hig
+ 964.500000n V_hig
+ 964.500001n V_hig
+ 964.600000n V_hig
+ 964.600001n V_hig
+ 964.700000n V_hig
+ 964.700001n V_hig
+ 964.800000n V_hig
+ 964.800001n V_hig
+ 964.900000n V_hig
+ 964.900001n V_hig
+ 965.000000n V_hig
+ 965.000001n V_low
+ 965.100000n V_low
+ 965.100001n V_low
+ 965.200000n V_low
+ 965.200001n V_low
+ 965.300000n V_low
+ 965.300001n V_low
+ 965.400000n V_low
+ 965.400001n V_low
+ 965.500000n V_low
+ 965.500001n V_low
+ 965.600000n V_low
+ 965.600001n V_low
+ 965.700000n V_low
+ 965.700001n V_low
+ 965.800000n V_low
+ 965.800001n V_low
+ 965.900000n V_low
+ 965.900001n V_low
+ 966.000000n V_low
+ 966.000001n V_hig
+ 966.100000n V_hig
+ 966.100001n V_hig
+ 966.200000n V_hig
+ 966.200001n V_hig
+ 966.300000n V_hig
+ 966.300001n V_hig
+ 966.400000n V_hig
+ 966.400001n V_hig
+ 966.500000n V_hig
+ 966.500001n V_hig
+ 966.600000n V_hig
+ 966.600001n V_hig
+ 966.700000n V_hig
+ 966.700001n V_hig
+ 966.800000n V_hig
+ 966.800001n V_hig
+ 966.900000n V_hig
+ 966.900001n V_hig
+ 967.000000n V_hig
+ 967.000001n V_low
+ 967.100000n V_low
+ 967.100001n V_low
+ 967.200000n V_low
+ 967.200001n V_low
+ 967.300000n V_low
+ 967.300001n V_low
+ 967.400000n V_low
+ 967.400001n V_low
+ 967.500000n V_low
+ 967.500001n V_low
+ 967.600000n V_low
+ 967.600001n V_low
+ 967.700000n V_low
+ 967.700001n V_low
+ 967.800000n V_low
+ 967.800001n V_low
+ 967.900000n V_low
+ 967.900001n V_low
+ 968.000000n V_low
+ 968.000001n V_low
+ 968.100000n V_low
+ 968.100001n V_low
+ 968.200000n V_low
+ 968.200001n V_low
+ 968.300000n V_low
+ 968.300001n V_low
+ 968.400000n V_low
+ 968.400001n V_low
+ 968.500000n V_low
+ 968.500001n V_low
+ 968.600000n V_low
+ 968.600001n V_low
+ 968.700000n V_low
+ 968.700001n V_low
+ 968.800000n V_low
+ 968.800001n V_low
+ 968.900000n V_low
+ 968.900001n V_low
+ 969.000000n V_low
+ 969.000001n V_hig
+ 969.100000n V_hig
+ 969.100001n V_hig
+ 969.200000n V_hig
+ 969.200001n V_hig
+ 969.300000n V_hig
+ 969.300001n V_hig
+ 969.400000n V_hig
+ 969.400001n V_hig
+ 969.500000n V_hig
+ 969.500001n V_hig
+ 969.600000n V_hig
+ 969.600001n V_hig
+ 969.700000n V_hig
+ 969.700001n V_hig
+ 969.800000n V_hig
+ 969.800001n V_hig
+ 969.900000n V_hig
+ 969.900001n V_hig
+ 970.000000n V_hig
+ 970.000001n V_low
+ 970.100000n V_low
+ 970.100001n V_low
+ 970.200000n V_low
+ 970.200001n V_low
+ 970.300000n V_low
+ 970.300001n V_low
+ 970.400000n V_low
+ 970.400001n V_low
+ 970.500000n V_low
+ 970.500001n V_low
+ 970.600000n V_low
+ 970.600001n V_low
+ 970.700000n V_low
+ 970.700001n V_low
+ 970.800000n V_low
+ 970.800001n V_low
+ 970.900000n V_low
+ 970.900001n V_low
+ 971.000000n V_low
+ 971.000001n V_hig
+ 971.100000n V_hig
+ 971.100001n V_hig
+ 971.200000n V_hig
+ 971.200001n V_hig
+ 971.300000n V_hig
+ 971.300001n V_hig
+ 971.400000n V_hig
+ 971.400001n V_hig
+ 971.500000n V_hig
+ 971.500001n V_hig
+ 971.600000n V_hig
+ 971.600001n V_hig
+ 971.700000n V_hig
+ 971.700001n V_hig
+ 971.800000n V_hig
+ 971.800001n V_hig
+ 971.900000n V_hig
+ 971.900001n V_hig
+ 972.000000n V_hig
+ 972.000001n V_hig
+ 972.100000n V_hig
+ 972.100001n V_hig
+ 972.200000n V_hig
+ 972.200001n V_hig
+ 972.300000n V_hig
+ 972.300001n V_hig
+ 972.400000n V_hig
+ 972.400001n V_hig
+ 972.500000n V_hig
+ 972.500001n V_hig
+ 972.600000n V_hig
+ 972.600001n V_hig
+ 972.700000n V_hig
+ 972.700001n V_hig
+ 972.800000n V_hig
+ 972.800001n V_hig
+ 972.900000n V_hig
+ 972.900001n V_hig
+ 973.000000n V_hig
+ 973.000001n V_low
+ 973.100000n V_low
+ 973.100001n V_low
+ 973.200000n V_low
+ 973.200001n V_low
+ 973.300000n V_low
+ 973.300001n V_low
+ 973.400000n V_low
+ 973.400001n V_low
+ 973.500000n V_low
+ 973.500001n V_low
+ 973.600000n V_low
+ 973.600001n V_low
+ 973.700000n V_low
+ 973.700001n V_low
+ 973.800000n V_low
+ 973.800001n V_low
+ 973.900000n V_low
+ 973.900001n V_low
+ 974.000000n V_low
+ 974.000001n V_hig
+ 974.100000n V_hig
+ 974.100001n V_hig
+ 974.200000n V_hig
+ 974.200001n V_hig
+ 974.300000n V_hig
+ 974.300001n V_hig
+ 974.400000n V_hig
+ 974.400001n V_hig
+ 974.500000n V_hig
+ 974.500001n V_hig
+ 974.600000n V_hig
+ 974.600001n V_hig
+ 974.700000n V_hig
+ 974.700001n V_hig
+ 974.800000n V_hig
+ 974.800001n V_hig
+ 974.900000n V_hig
+ 974.900001n V_hig
+ 975.000000n V_hig
+ 975.000001n V_low
+ 975.100000n V_low
+ 975.100001n V_low
+ 975.200000n V_low
+ 975.200001n V_low
+ 975.300000n V_low
+ 975.300001n V_low
+ 975.400000n V_low
+ 975.400001n V_low
+ 975.500000n V_low
+ 975.500001n V_low
+ 975.600000n V_low
+ 975.600001n V_low
+ 975.700000n V_low
+ 975.700001n V_low
+ 975.800000n V_low
+ 975.800001n V_low
+ 975.900000n V_low
+ 975.900001n V_low
+ 976.000000n V_low
+ 976.000001n V_low
+ 976.100000n V_low
+ 976.100001n V_low
+ 976.200000n V_low
+ 976.200001n V_low
+ 976.300000n V_low
+ 976.300001n V_low
+ 976.400000n V_low
+ 976.400001n V_low
+ 976.500000n V_low
+ 976.500001n V_low
+ 976.600000n V_low
+ 976.600001n V_low
+ 976.700000n V_low
+ 976.700001n V_low
+ 976.800000n V_low
+ 976.800001n V_low
+ 976.900000n V_low
+ 976.900001n V_low
+ 977.000000n V_low
+ 977.000001n V_hig
+ 977.100000n V_hig
+ 977.100001n V_hig
+ 977.200000n V_hig
+ 977.200001n V_hig
+ 977.300000n V_hig
+ 977.300001n V_hig
+ 977.400000n V_hig
+ 977.400001n V_hig
+ 977.500000n V_hig
+ 977.500001n V_hig
+ 977.600000n V_hig
+ 977.600001n V_hig
+ 977.700000n V_hig
+ 977.700001n V_hig
+ 977.800000n V_hig
+ 977.800001n V_hig
+ 977.900000n V_hig
+ 977.900001n V_hig
+ 978.000000n V_hig
+ 978.000001n V_hig
+ 978.100000n V_hig
+ 978.100001n V_hig
+ 978.200000n V_hig
+ 978.200001n V_hig
+ 978.300000n V_hig
+ 978.300001n V_hig
+ 978.400000n V_hig
+ 978.400001n V_hig
+ 978.500000n V_hig
+ 978.500001n V_hig
+ 978.600000n V_hig
+ 978.600001n V_hig
+ 978.700000n V_hig
+ 978.700001n V_hig
+ 978.800000n V_hig
+ 978.800001n V_hig
+ 978.900000n V_hig
+ 978.900001n V_hig
+ 979.000000n V_hig
+ 979.000001n V_low
+ 979.100000n V_low
+ 979.100001n V_low
+ 979.200000n V_low
+ 979.200001n V_low
+ 979.300000n V_low
+ 979.300001n V_low
+ 979.400000n V_low
+ 979.400001n V_low
+ 979.500000n V_low
+ 979.500001n V_low
+ 979.600000n V_low
+ 979.600001n V_low
+ 979.700000n V_low
+ 979.700001n V_low
+ 979.800000n V_low
+ 979.800001n V_low
+ 979.900000n V_low
+ 979.900001n V_low
+ 980.000000n V_low
+ 980.000001n V_hig
+ 980.100000n V_hig
+ 980.100001n V_hig
+ 980.200000n V_hig
+ 980.200001n V_hig
+ 980.300000n V_hig
+ 980.300001n V_hig
+ 980.400000n V_hig
+ 980.400001n V_hig
+ 980.500000n V_hig
+ 980.500001n V_hig
+ 980.600000n V_hig
+ 980.600001n V_hig
+ 980.700000n V_hig
+ 980.700001n V_hig
+ 980.800000n V_hig
+ 980.800001n V_hig
+ 980.900000n V_hig
+ 980.900001n V_hig
+ 981.000000n V_hig
+ 981.000001n V_hig
+ 981.100000n V_hig
+ 981.100001n V_hig
+ 981.200000n V_hig
+ 981.200001n V_hig
+ 981.300000n V_hig
+ 981.300001n V_hig
+ 981.400000n V_hig
+ 981.400001n V_hig
+ 981.500000n V_hig
+ 981.500001n V_hig
+ 981.600000n V_hig
+ 981.600001n V_hig
+ 981.700000n V_hig
+ 981.700001n V_hig
+ 981.800000n V_hig
+ 981.800001n V_hig
+ 981.900000n V_hig
+ 981.900001n V_hig
+ 982.000000n V_hig
+ 982.000001n V_low
+ 982.100000n V_low
+ 982.100001n V_low
+ 982.200000n V_low
+ 982.200001n V_low
+ 982.300000n V_low
+ 982.300001n V_low
+ 982.400000n V_low
+ 982.400001n V_low
+ 982.500000n V_low
+ 982.500001n V_low
+ 982.600000n V_low
+ 982.600001n V_low
+ 982.700000n V_low
+ 982.700001n V_low
+ 982.800000n V_low
+ 982.800001n V_low
+ 982.900000n V_low
+ 982.900001n V_low
+ 983.000000n V_low
+ 983.000001n V_hig
+ 983.100000n V_hig
+ 983.100001n V_hig
+ 983.200000n V_hig
+ 983.200001n V_hig
+ 983.300000n V_hig
+ 983.300001n V_hig
+ 983.400000n V_hig
+ 983.400001n V_hig
+ 983.500000n V_hig
+ 983.500001n V_hig
+ 983.600000n V_hig
+ 983.600001n V_hig
+ 983.700000n V_hig
+ 983.700001n V_hig
+ 983.800000n V_hig
+ 983.800001n V_hig
+ 983.900000n V_hig
+ 983.900001n V_hig
+ 984.000000n V_hig
+ 984.000001n V_low
+ 984.100000n V_low
+ 984.100001n V_low
+ 984.200000n V_low
+ 984.200001n V_low
+ 984.300000n V_low
+ 984.300001n V_low
+ 984.400000n V_low
+ 984.400001n V_low
+ 984.500000n V_low
+ 984.500001n V_low
+ 984.600000n V_low
+ 984.600001n V_low
+ 984.700000n V_low
+ 984.700001n V_low
+ 984.800000n V_low
+ 984.800001n V_low
+ 984.900000n V_low
+ 984.900001n V_low
+ 985.000000n V_low
+ 985.000001n V_low
+ 985.100000n V_low
+ 985.100001n V_low
+ 985.200000n V_low
+ 985.200001n V_low
+ 985.300000n V_low
+ 985.300001n V_low
+ 985.400000n V_low
+ 985.400001n V_low
+ 985.500000n V_low
+ 985.500001n V_low
+ 985.600000n V_low
+ 985.600001n V_low
+ 985.700000n V_low
+ 985.700001n V_low
+ 985.800000n V_low
+ 985.800001n V_low
+ 985.900000n V_low
+ 985.900001n V_low
+ 986.000000n V_low
+ 986.000001n V_low
+ 986.100000n V_low
+ 986.100001n V_low
+ 986.200000n V_low
+ 986.200001n V_low
+ 986.300000n V_low
+ 986.300001n V_low
+ 986.400000n V_low
+ 986.400001n V_low
+ 986.500000n V_low
+ 986.500001n V_low
+ 986.600000n V_low
+ 986.600001n V_low
+ 986.700000n V_low
+ 986.700001n V_low
+ 986.800000n V_low
+ 986.800001n V_low
+ 986.900000n V_low
+ 986.900001n V_low
+ 987.000000n V_low
+ 987.000001n V_hig
+ 987.100000n V_hig
+ 987.100001n V_hig
+ 987.200000n V_hig
+ 987.200001n V_hig
+ 987.300000n V_hig
+ 987.300001n V_hig
+ 987.400000n V_hig
+ 987.400001n V_hig
+ 987.500000n V_hig
+ 987.500001n V_hig
+ 987.600000n V_hig
+ 987.600001n V_hig
+ 987.700000n V_hig
+ 987.700001n V_hig
+ 987.800000n V_hig
+ 987.800001n V_hig
+ 987.900000n V_hig
+ 987.900001n V_hig
+ 988.000000n V_hig
+ 988.000001n V_hig
+ 988.100000n V_hig
+ 988.100001n V_hig
+ 988.200000n V_hig
+ 988.200001n V_hig
+ 988.300000n V_hig
+ 988.300001n V_hig
+ 988.400000n V_hig
+ 988.400001n V_hig
+ 988.500000n V_hig
+ 988.500001n V_hig
+ 988.600000n V_hig
+ 988.600001n V_hig
+ 988.700000n V_hig
+ 988.700001n V_hig
+ 988.800000n V_hig
+ 988.800001n V_hig
+ 988.900000n V_hig
+ 988.900001n V_hig
+ 989.000000n V_hig
+ 989.000001n V_hig
+ 989.100000n V_hig
+ 989.100001n V_hig
+ 989.200000n V_hig
+ 989.200001n V_hig
+ 989.300000n V_hig
+ 989.300001n V_hig
+ 989.400000n V_hig
+ 989.400001n V_hig
+ 989.500000n V_hig
+ 989.500001n V_hig
+ 989.600000n V_hig
+ 989.600001n V_hig
+ 989.700000n V_hig
+ 989.700001n V_hig
+ 989.800000n V_hig
+ 989.800001n V_hig
+ 989.900000n V_hig
+ 989.900001n V_hig
+ 990.000000n V_hig
+ 990.000001n V_hig
+ 990.100000n V_hig
+ 990.100001n V_hig
+ 990.200000n V_hig
+ 990.200001n V_hig
+ 990.300000n V_hig
+ 990.300001n V_hig
+ 990.400000n V_hig
+ 990.400001n V_hig
+ 990.500000n V_hig
+ 990.500001n V_hig
+ 990.600000n V_hig
+ 990.600001n V_hig
+ 990.700000n V_hig
+ 990.700001n V_hig
+ 990.800000n V_hig
+ 990.800001n V_hig
+ 990.900000n V_hig
+ 990.900001n V_hig
+ 991.000000n V_hig
+ 991.000001n V_hig
+ 991.100000n V_hig
+ 991.100001n V_hig
+ 991.200000n V_hig
+ 991.200001n V_hig
+ 991.300000n V_hig
+ 991.300001n V_hig
+ 991.400000n V_hig
+ 991.400001n V_hig
+ 991.500000n V_hig
+ 991.500001n V_hig
+ 991.600000n V_hig
+ 991.600001n V_hig
+ 991.700000n V_hig
+ 991.700001n V_hig
+ 991.800000n V_hig
+ 991.800001n V_hig
+ 991.900000n V_hig
+ 991.900001n V_hig
+ 992.000000n V_hig
+ 992.000001n V_low
+ 992.100000n V_low
+ 992.100001n V_low
+ 992.200000n V_low
+ 992.200001n V_low
+ 992.300000n V_low
+ 992.300001n V_low
+ 992.400000n V_low
+ 992.400001n V_low
+ 992.500000n V_low
+ 992.500001n V_low
+ 992.600000n V_low
+ 992.600001n V_low
+ 992.700000n V_low
+ 992.700001n V_low
+ 992.800000n V_low
+ 992.800001n V_low
+ 992.900000n V_low
+ 992.900001n V_low
+ 993.000000n V_low
+ 993.000001n V_hig
+ 993.100000n V_hig
+ 993.100001n V_hig
+ 993.200000n V_hig
+ 993.200001n V_hig
+ 993.300000n V_hig
+ 993.300001n V_hig
+ 993.400000n V_hig
+ 993.400001n V_hig
+ 993.500000n V_hig
+ 993.500001n V_hig
+ 993.600000n V_hig
+ 993.600001n V_hig
+ 993.700000n V_hig
+ 993.700001n V_hig
+ 993.800000n V_hig
+ 993.800001n V_hig
+ 993.900000n V_hig
+ 993.900001n V_hig
+ 994.000000n V_hig
+ 994.000001n V_low
+ 994.100000n V_low
+ 994.100001n V_low
+ 994.200000n V_low
+ 994.200001n V_low
+ 994.300000n V_low
+ 994.300001n V_low
+ 994.400000n V_low
+ 994.400001n V_low
+ 994.500000n V_low
+ 994.500001n V_low
+ 994.600000n V_low
+ 994.600001n V_low
+ 994.700000n V_low
+ 994.700001n V_low
+ 994.800000n V_low
+ 994.800001n V_low
+ 994.900000n V_low
+ 994.900001n V_low
+ 995.000000n V_low
+ 995.000001n V_low
+ 995.100000n V_low
+ 995.100001n V_low
+ 995.200000n V_low
+ 995.200001n V_low
+ 995.300000n V_low
+ 995.300001n V_low
+ 995.400000n V_low
+ 995.400001n V_low
+ 995.500000n V_low
+ 995.500001n V_low
+ 995.600000n V_low
+ 995.600001n V_low
+ 995.700000n V_low
+ 995.700001n V_low
+ 995.800000n V_low
+ 995.800001n V_low
+ 995.900000n V_low
+ 995.900001n V_low
+ 996.000000n V_low
+ 996.000001n V_low
+ 996.100000n V_low
+ 996.100001n V_low
+ 996.200000n V_low
+ 996.200001n V_low
+ 996.300000n V_low
+ 996.300001n V_low
+ 996.400000n V_low
+ 996.400001n V_low
+ 996.500000n V_low
+ 996.500001n V_low
+ 996.600000n V_low
+ 996.600001n V_low
+ 996.700000n V_low
+ 996.700001n V_low
+ 996.800000n V_low
+ 996.800001n V_low
+ 996.900000n V_low
+ 996.900001n V_low
+ 997.000000n V_low
+ 997.000001n V_low
+ 997.100000n V_low
+ 997.100001n V_low
+ 997.200000n V_low
+ 997.200001n V_low
+ 997.300000n V_low
+ 997.300001n V_low
+ 997.400000n V_low
+ 997.400001n V_low
+ 997.500000n V_low
+ 997.500001n V_low
+ 997.600000n V_low
+ 997.600001n V_low
+ 997.700000n V_low
+ 997.700001n V_low
+ 997.800000n V_low
+ 997.800001n V_low
+ 997.900000n V_low
+ 997.900001n V_low
+ 998.000000n V_low
+ 998.000001n V_low
+ 998.100000n V_low
+ 998.100001n V_low
+ 998.200000n V_low
+ 998.200001n V_low
+ 998.300000n V_low
+ 998.300001n V_low
+ 998.400000n V_low
+ 998.400001n V_low
+ 998.500000n V_low
+ 998.500001n V_low
+ 998.600000n V_low
+ 998.600001n V_low
+ 998.700000n V_low
+ 998.700001n V_low
+ 998.800000n V_low
+ 998.800001n V_low
+ 998.900000n V_low
+ 998.900001n V_low
+ 999.000000n V_low
+ 999.000001n V_hig
+ 999.100000n V_hig
+ 999.100001n V_hig
+ 999.200000n V_hig
+ 999.200001n V_hig
+ 999.300000n V_hig
+ 999.300001n V_hig
+ 999.400000n V_hig
+ 999.400001n V_hig
+ 999.500000n V_hig
+ 999.500001n V_hig
+ 999.600000n V_hig
+ 999.600001n V_hig
+ 999.700000n V_hig
+ 999.700001n V_hig
+ 999.800000n V_hig
+ 999.800001n V_hig
+ 999.900000n V_hig
+ 999.900001n V_hig
+ 1000.000000n V_hig
+ 
v2 b1 0 PWL
+ 0.000001n V_low
+ 0.100000n V_low
+ 0.100001n V_low
+ 0.200000n V_low
+ 0.200001n V_low
+ 0.300000n V_low
+ 0.300001n V_low
+ 0.400000n V_low
+ 0.400001n V_low
+ 0.500000n V_low
+ 0.500001n V_low
+ 0.600000n V_low
+ 0.600001n V_low
+ 0.700000n V_low
+ 0.700001n V_low
+ 0.800000n V_low
+ 0.800001n V_low
+ 0.900000n V_low
+ 0.900001n V_low
+ 1.000000n V_low
+ 1.000001n V_low
+ 1.100000n V_low
+ 1.100001n V_low
+ 1.200000n V_low
+ 1.200001n V_low
+ 1.300000n V_low
+ 1.300001n V_low
+ 1.400000n V_low
+ 1.400001n V_low
+ 1.500000n V_low
+ 1.500001n V_low
+ 1.600000n V_low
+ 1.600001n V_low
+ 1.700000n V_low
+ 1.700001n V_low
+ 1.800000n V_low
+ 1.800001n V_low
+ 1.900000n V_low
+ 1.900001n V_low
+ 2.000000n V_low
+ 2.000001n V_low
+ 2.100000n V_low
+ 2.100001n V_low
+ 2.200000n V_low
+ 2.200001n V_low
+ 2.300000n V_low
+ 2.300001n V_low
+ 2.400000n V_low
+ 2.400001n V_low
+ 2.500000n V_low
+ 2.500001n V_low
+ 2.600000n V_low
+ 2.600001n V_low
+ 2.700000n V_low
+ 2.700001n V_low
+ 2.800000n V_low
+ 2.800001n V_low
+ 2.900000n V_low
+ 2.900001n V_low
+ 3.000000n V_low
+ 3.000001n V_low
+ 3.100000n V_low
+ 3.100001n V_low
+ 3.200000n V_low
+ 3.200001n V_low
+ 3.300000n V_low
+ 3.300001n V_low
+ 3.400000n V_low
+ 3.400001n V_low
+ 3.500000n V_low
+ 3.500001n V_low
+ 3.600000n V_low
+ 3.600001n V_low
+ 3.700000n V_low
+ 3.700001n V_low
+ 3.800000n V_low
+ 3.800001n V_low
+ 3.900000n V_low
+ 3.900001n V_low
+ 4.000000n V_low
+ 4.000001n V_hig
+ 4.100000n V_hig
+ 4.100001n V_hig
+ 4.200000n V_hig
+ 4.200001n V_hig
+ 4.300000n V_hig
+ 4.300001n V_hig
+ 4.400000n V_hig
+ 4.400001n V_hig
+ 4.500000n V_hig
+ 4.500001n V_hig
+ 4.600000n V_hig
+ 4.600001n V_hig
+ 4.700000n V_hig
+ 4.700001n V_hig
+ 4.800000n V_hig
+ 4.800001n V_hig
+ 4.900000n V_hig
+ 4.900001n V_hig
+ 5.000000n V_hig
+ 5.000001n V_hig
+ 5.100000n V_hig
+ 5.100001n V_hig
+ 5.200000n V_hig
+ 5.200001n V_hig
+ 5.300000n V_hig
+ 5.300001n V_hig
+ 5.400000n V_hig
+ 5.400001n V_hig
+ 5.500000n V_hig
+ 5.500001n V_hig
+ 5.600000n V_hig
+ 5.600001n V_hig
+ 5.700000n V_hig
+ 5.700001n V_hig
+ 5.800000n V_hig
+ 5.800001n V_hig
+ 5.900000n V_hig
+ 5.900001n V_hig
+ 6.000000n V_hig
+ 6.000001n V_hig
+ 6.100000n V_hig
+ 6.100001n V_hig
+ 6.200000n V_hig
+ 6.200001n V_hig
+ 6.300000n V_hig
+ 6.300001n V_hig
+ 6.400000n V_hig
+ 6.400001n V_hig
+ 6.500000n V_hig
+ 6.500001n V_hig
+ 6.600000n V_hig
+ 6.600001n V_hig
+ 6.700000n V_hig
+ 6.700001n V_hig
+ 6.800000n V_hig
+ 6.800001n V_hig
+ 6.900000n V_hig
+ 6.900001n V_hig
+ 7.000000n V_hig
+ 7.000001n V_hig
+ 7.100000n V_hig
+ 7.100001n V_hig
+ 7.200000n V_hig
+ 7.200001n V_hig
+ 7.300000n V_hig
+ 7.300001n V_hig
+ 7.400000n V_hig
+ 7.400001n V_hig
+ 7.500000n V_hig
+ 7.500001n V_hig
+ 7.600000n V_hig
+ 7.600001n V_hig
+ 7.700000n V_hig
+ 7.700001n V_hig
+ 7.800000n V_hig
+ 7.800001n V_hig
+ 7.900000n V_hig
+ 7.900001n V_hig
+ 8.000000n V_hig
+ 8.000001n V_hig
+ 8.100000n V_hig
+ 8.100001n V_hig
+ 8.200000n V_hig
+ 8.200001n V_hig
+ 8.300000n V_hig
+ 8.300001n V_hig
+ 8.400000n V_hig
+ 8.400001n V_hig
+ 8.500000n V_hig
+ 8.500001n V_hig
+ 8.600000n V_hig
+ 8.600001n V_hig
+ 8.700000n V_hig
+ 8.700001n V_hig
+ 8.800000n V_hig
+ 8.800001n V_hig
+ 8.900000n V_hig
+ 8.900001n V_hig
+ 9.000000n V_hig
+ 9.000001n V_hig
+ 9.100000n V_hig
+ 9.100001n V_hig
+ 9.200000n V_hig
+ 9.200001n V_hig
+ 9.300000n V_hig
+ 9.300001n V_hig
+ 9.400000n V_hig
+ 9.400001n V_hig
+ 9.500000n V_hig
+ 9.500001n V_hig
+ 9.600000n V_hig
+ 9.600001n V_hig
+ 9.700000n V_hig
+ 9.700001n V_hig
+ 9.800000n V_hig
+ 9.800001n V_hig
+ 9.900000n V_hig
+ 9.900001n V_hig
+ 10.000000n V_hig
+ 10.000001n V_low
+ 10.100000n V_low
+ 10.100001n V_low
+ 10.200000n V_low
+ 10.200001n V_low
+ 10.300000n V_low
+ 10.300001n V_low
+ 10.400000n V_low
+ 10.400001n V_low
+ 10.500000n V_low
+ 10.500001n V_low
+ 10.600000n V_low
+ 10.600001n V_low
+ 10.700000n V_low
+ 10.700001n V_low
+ 10.800000n V_low
+ 10.800001n V_low
+ 10.900000n V_low
+ 10.900001n V_low
+ 11.000000n V_low
+ 11.000001n V_hig
+ 11.100000n V_hig
+ 11.100001n V_hig
+ 11.200000n V_hig
+ 11.200001n V_hig
+ 11.300000n V_hig
+ 11.300001n V_hig
+ 11.400000n V_hig
+ 11.400001n V_hig
+ 11.500000n V_hig
+ 11.500001n V_hig
+ 11.600000n V_hig
+ 11.600001n V_hig
+ 11.700000n V_hig
+ 11.700001n V_hig
+ 11.800000n V_hig
+ 11.800001n V_hig
+ 11.900000n V_hig
+ 11.900001n V_hig
+ 12.000000n V_hig
+ 12.000001n V_hig
+ 12.100000n V_hig
+ 12.100001n V_hig
+ 12.200000n V_hig
+ 12.200001n V_hig
+ 12.300000n V_hig
+ 12.300001n V_hig
+ 12.400000n V_hig
+ 12.400001n V_hig
+ 12.500000n V_hig
+ 12.500001n V_hig
+ 12.600000n V_hig
+ 12.600001n V_hig
+ 12.700000n V_hig
+ 12.700001n V_hig
+ 12.800000n V_hig
+ 12.800001n V_hig
+ 12.900000n V_hig
+ 12.900001n V_hig
+ 13.000000n V_hig
+ 13.000001n V_low
+ 13.100000n V_low
+ 13.100001n V_low
+ 13.200000n V_low
+ 13.200001n V_low
+ 13.300000n V_low
+ 13.300001n V_low
+ 13.400000n V_low
+ 13.400001n V_low
+ 13.500000n V_low
+ 13.500001n V_low
+ 13.600000n V_low
+ 13.600001n V_low
+ 13.700000n V_low
+ 13.700001n V_low
+ 13.800000n V_low
+ 13.800001n V_low
+ 13.900000n V_low
+ 13.900001n V_low
+ 14.000000n V_low
+ 14.000001n V_hig
+ 14.100000n V_hig
+ 14.100001n V_hig
+ 14.200000n V_hig
+ 14.200001n V_hig
+ 14.300000n V_hig
+ 14.300001n V_hig
+ 14.400000n V_hig
+ 14.400001n V_hig
+ 14.500000n V_hig
+ 14.500001n V_hig
+ 14.600000n V_hig
+ 14.600001n V_hig
+ 14.700000n V_hig
+ 14.700001n V_hig
+ 14.800000n V_hig
+ 14.800001n V_hig
+ 14.900000n V_hig
+ 14.900001n V_hig
+ 15.000000n V_hig
+ 15.000001n V_low
+ 15.100000n V_low
+ 15.100001n V_low
+ 15.200000n V_low
+ 15.200001n V_low
+ 15.300000n V_low
+ 15.300001n V_low
+ 15.400000n V_low
+ 15.400001n V_low
+ 15.500000n V_low
+ 15.500001n V_low
+ 15.600000n V_low
+ 15.600001n V_low
+ 15.700000n V_low
+ 15.700001n V_low
+ 15.800000n V_low
+ 15.800001n V_low
+ 15.900000n V_low
+ 15.900001n V_low
+ 16.000000n V_low
+ 16.000001n V_hig
+ 16.100000n V_hig
+ 16.100001n V_hig
+ 16.200000n V_hig
+ 16.200001n V_hig
+ 16.300000n V_hig
+ 16.300001n V_hig
+ 16.400000n V_hig
+ 16.400001n V_hig
+ 16.500000n V_hig
+ 16.500001n V_hig
+ 16.600000n V_hig
+ 16.600001n V_hig
+ 16.700000n V_hig
+ 16.700001n V_hig
+ 16.800000n V_hig
+ 16.800001n V_hig
+ 16.900000n V_hig
+ 16.900001n V_hig
+ 17.000000n V_hig
+ 17.000001n V_hig
+ 17.100000n V_hig
+ 17.100001n V_hig
+ 17.200000n V_hig
+ 17.200001n V_hig
+ 17.300000n V_hig
+ 17.300001n V_hig
+ 17.400000n V_hig
+ 17.400001n V_hig
+ 17.500000n V_hig
+ 17.500001n V_hig
+ 17.600000n V_hig
+ 17.600001n V_hig
+ 17.700000n V_hig
+ 17.700001n V_hig
+ 17.800000n V_hig
+ 17.800001n V_hig
+ 17.900000n V_hig
+ 17.900001n V_hig
+ 18.000000n V_hig
+ 18.000001n V_low
+ 18.100000n V_low
+ 18.100001n V_low
+ 18.200000n V_low
+ 18.200001n V_low
+ 18.300000n V_low
+ 18.300001n V_low
+ 18.400000n V_low
+ 18.400001n V_low
+ 18.500000n V_low
+ 18.500001n V_low
+ 18.600000n V_low
+ 18.600001n V_low
+ 18.700000n V_low
+ 18.700001n V_low
+ 18.800000n V_low
+ 18.800001n V_low
+ 18.900000n V_low
+ 18.900001n V_low
+ 19.000000n V_low
+ 19.000001n V_low
+ 19.100000n V_low
+ 19.100001n V_low
+ 19.200000n V_low
+ 19.200001n V_low
+ 19.300000n V_low
+ 19.300001n V_low
+ 19.400000n V_low
+ 19.400001n V_low
+ 19.500000n V_low
+ 19.500001n V_low
+ 19.600000n V_low
+ 19.600001n V_low
+ 19.700000n V_low
+ 19.700001n V_low
+ 19.800000n V_low
+ 19.800001n V_low
+ 19.900000n V_low
+ 19.900001n V_low
+ 20.000000n V_low
+ 20.000001n V_hig
+ 20.100000n V_hig
+ 20.100001n V_hig
+ 20.200000n V_hig
+ 20.200001n V_hig
+ 20.300000n V_hig
+ 20.300001n V_hig
+ 20.400000n V_hig
+ 20.400001n V_hig
+ 20.500000n V_hig
+ 20.500001n V_hig
+ 20.600000n V_hig
+ 20.600001n V_hig
+ 20.700000n V_hig
+ 20.700001n V_hig
+ 20.800000n V_hig
+ 20.800001n V_hig
+ 20.900000n V_hig
+ 20.900001n V_hig
+ 21.000000n V_hig
+ 21.000001n V_hig
+ 21.100000n V_hig
+ 21.100001n V_hig
+ 21.200000n V_hig
+ 21.200001n V_hig
+ 21.300000n V_hig
+ 21.300001n V_hig
+ 21.400000n V_hig
+ 21.400001n V_hig
+ 21.500000n V_hig
+ 21.500001n V_hig
+ 21.600000n V_hig
+ 21.600001n V_hig
+ 21.700000n V_hig
+ 21.700001n V_hig
+ 21.800000n V_hig
+ 21.800001n V_hig
+ 21.900000n V_hig
+ 21.900001n V_hig
+ 22.000000n V_hig
+ 22.000001n V_hig
+ 22.100000n V_hig
+ 22.100001n V_hig
+ 22.200000n V_hig
+ 22.200001n V_hig
+ 22.300000n V_hig
+ 22.300001n V_hig
+ 22.400000n V_hig
+ 22.400001n V_hig
+ 22.500000n V_hig
+ 22.500001n V_hig
+ 22.600000n V_hig
+ 22.600001n V_hig
+ 22.700000n V_hig
+ 22.700001n V_hig
+ 22.800000n V_hig
+ 22.800001n V_hig
+ 22.900000n V_hig
+ 22.900001n V_hig
+ 23.000000n V_hig
+ 23.000001n V_hig
+ 23.100000n V_hig
+ 23.100001n V_hig
+ 23.200000n V_hig
+ 23.200001n V_hig
+ 23.300000n V_hig
+ 23.300001n V_hig
+ 23.400000n V_hig
+ 23.400001n V_hig
+ 23.500000n V_hig
+ 23.500001n V_hig
+ 23.600000n V_hig
+ 23.600001n V_hig
+ 23.700000n V_hig
+ 23.700001n V_hig
+ 23.800000n V_hig
+ 23.800001n V_hig
+ 23.900000n V_hig
+ 23.900001n V_hig
+ 24.000000n V_hig
+ 24.000001n V_low
+ 24.100000n V_low
+ 24.100001n V_low
+ 24.200000n V_low
+ 24.200001n V_low
+ 24.300000n V_low
+ 24.300001n V_low
+ 24.400000n V_low
+ 24.400001n V_low
+ 24.500000n V_low
+ 24.500001n V_low
+ 24.600000n V_low
+ 24.600001n V_low
+ 24.700000n V_low
+ 24.700001n V_low
+ 24.800000n V_low
+ 24.800001n V_low
+ 24.900000n V_low
+ 24.900001n V_low
+ 25.000000n V_low
+ 25.000001n V_low
+ 25.100000n V_low
+ 25.100001n V_low
+ 25.200000n V_low
+ 25.200001n V_low
+ 25.300000n V_low
+ 25.300001n V_low
+ 25.400000n V_low
+ 25.400001n V_low
+ 25.500000n V_low
+ 25.500001n V_low
+ 25.600000n V_low
+ 25.600001n V_low
+ 25.700000n V_low
+ 25.700001n V_low
+ 25.800000n V_low
+ 25.800001n V_low
+ 25.900000n V_low
+ 25.900001n V_low
+ 26.000000n V_low
+ 26.000001n V_hig
+ 26.100000n V_hig
+ 26.100001n V_hig
+ 26.200000n V_hig
+ 26.200001n V_hig
+ 26.300000n V_hig
+ 26.300001n V_hig
+ 26.400000n V_hig
+ 26.400001n V_hig
+ 26.500000n V_hig
+ 26.500001n V_hig
+ 26.600000n V_hig
+ 26.600001n V_hig
+ 26.700000n V_hig
+ 26.700001n V_hig
+ 26.800000n V_hig
+ 26.800001n V_hig
+ 26.900000n V_hig
+ 26.900001n V_hig
+ 27.000000n V_hig
+ 27.000001n V_hig
+ 27.100000n V_hig
+ 27.100001n V_hig
+ 27.200000n V_hig
+ 27.200001n V_hig
+ 27.300000n V_hig
+ 27.300001n V_hig
+ 27.400000n V_hig
+ 27.400001n V_hig
+ 27.500000n V_hig
+ 27.500001n V_hig
+ 27.600000n V_hig
+ 27.600001n V_hig
+ 27.700000n V_hig
+ 27.700001n V_hig
+ 27.800000n V_hig
+ 27.800001n V_hig
+ 27.900000n V_hig
+ 27.900001n V_hig
+ 28.000000n V_hig
+ 28.000001n V_hig
+ 28.100000n V_hig
+ 28.100001n V_hig
+ 28.200000n V_hig
+ 28.200001n V_hig
+ 28.300000n V_hig
+ 28.300001n V_hig
+ 28.400000n V_hig
+ 28.400001n V_hig
+ 28.500000n V_hig
+ 28.500001n V_hig
+ 28.600000n V_hig
+ 28.600001n V_hig
+ 28.700000n V_hig
+ 28.700001n V_hig
+ 28.800000n V_hig
+ 28.800001n V_hig
+ 28.900000n V_hig
+ 28.900001n V_hig
+ 29.000000n V_hig
+ 29.000001n V_low
+ 29.100000n V_low
+ 29.100001n V_low
+ 29.200000n V_low
+ 29.200001n V_low
+ 29.300000n V_low
+ 29.300001n V_low
+ 29.400000n V_low
+ 29.400001n V_low
+ 29.500000n V_low
+ 29.500001n V_low
+ 29.600000n V_low
+ 29.600001n V_low
+ 29.700000n V_low
+ 29.700001n V_low
+ 29.800000n V_low
+ 29.800001n V_low
+ 29.900000n V_low
+ 29.900001n V_low
+ 30.000000n V_low
+ 30.000001n V_low
+ 30.100000n V_low
+ 30.100001n V_low
+ 30.200000n V_low
+ 30.200001n V_low
+ 30.300000n V_low
+ 30.300001n V_low
+ 30.400000n V_low
+ 30.400001n V_low
+ 30.500000n V_low
+ 30.500001n V_low
+ 30.600000n V_low
+ 30.600001n V_low
+ 30.700000n V_low
+ 30.700001n V_low
+ 30.800000n V_low
+ 30.800001n V_low
+ 30.900000n V_low
+ 30.900001n V_low
+ 31.000000n V_low
+ 31.000001n V_low
+ 31.100000n V_low
+ 31.100001n V_low
+ 31.200000n V_low
+ 31.200001n V_low
+ 31.300000n V_low
+ 31.300001n V_low
+ 31.400000n V_low
+ 31.400001n V_low
+ 31.500000n V_low
+ 31.500001n V_low
+ 31.600000n V_low
+ 31.600001n V_low
+ 31.700000n V_low
+ 31.700001n V_low
+ 31.800000n V_low
+ 31.800001n V_low
+ 31.900000n V_low
+ 31.900001n V_low
+ 32.000000n V_low
+ 32.000001n V_low
+ 32.100000n V_low
+ 32.100001n V_low
+ 32.200000n V_low
+ 32.200001n V_low
+ 32.300000n V_low
+ 32.300001n V_low
+ 32.400000n V_low
+ 32.400001n V_low
+ 32.500000n V_low
+ 32.500001n V_low
+ 32.600000n V_low
+ 32.600001n V_low
+ 32.700000n V_low
+ 32.700001n V_low
+ 32.800000n V_low
+ 32.800001n V_low
+ 32.900000n V_low
+ 32.900001n V_low
+ 33.000000n V_low
+ 33.000001n V_low
+ 33.100000n V_low
+ 33.100001n V_low
+ 33.200000n V_low
+ 33.200001n V_low
+ 33.300000n V_low
+ 33.300001n V_low
+ 33.400000n V_low
+ 33.400001n V_low
+ 33.500000n V_low
+ 33.500001n V_low
+ 33.600000n V_low
+ 33.600001n V_low
+ 33.700000n V_low
+ 33.700001n V_low
+ 33.800000n V_low
+ 33.800001n V_low
+ 33.900000n V_low
+ 33.900001n V_low
+ 34.000000n V_low
+ 34.000001n V_hig
+ 34.100000n V_hig
+ 34.100001n V_hig
+ 34.200000n V_hig
+ 34.200001n V_hig
+ 34.300000n V_hig
+ 34.300001n V_hig
+ 34.400000n V_hig
+ 34.400001n V_hig
+ 34.500000n V_hig
+ 34.500001n V_hig
+ 34.600000n V_hig
+ 34.600001n V_hig
+ 34.700000n V_hig
+ 34.700001n V_hig
+ 34.800000n V_hig
+ 34.800001n V_hig
+ 34.900000n V_hig
+ 34.900001n V_hig
+ 35.000000n V_hig
+ 35.000001n V_low
+ 35.100000n V_low
+ 35.100001n V_low
+ 35.200000n V_low
+ 35.200001n V_low
+ 35.300000n V_low
+ 35.300001n V_low
+ 35.400000n V_low
+ 35.400001n V_low
+ 35.500000n V_low
+ 35.500001n V_low
+ 35.600000n V_low
+ 35.600001n V_low
+ 35.700000n V_low
+ 35.700001n V_low
+ 35.800000n V_low
+ 35.800001n V_low
+ 35.900000n V_low
+ 35.900001n V_low
+ 36.000000n V_low
+ 36.000001n V_low
+ 36.100000n V_low
+ 36.100001n V_low
+ 36.200000n V_low
+ 36.200001n V_low
+ 36.300000n V_low
+ 36.300001n V_low
+ 36.400000n V_low
+ 36.400001n V_low
+ 36.500000n V_low
+ 36.500001n V_low
+ 36.600000n V_low
+ 36.600001n V_low
+ 36.700000n V_low
+ 36.700001n V_low
+ 36.800000n V_low
+ 36.800001n V_low
+ 36.900000n V_low
+ 36.900001n V_low
+ 37.000000n V_low
+ 37.000001n V_hig
+ 37.100000n V_hig
+ 37.100001n V_hig
+ 37.200000n V_hig
+ 37.200001n V_hig
+ 37.300000n V_hig
+ 37.300001n V_hig
+ 37.400000n V_hig
+ 37.400001n V_hig
+ 37.500000n V_hig
+ 37.500001n V_hig
+ 37.600000n V_hig
+ 37.600001n V_hig
+ 37.700000n V_hig
+ 37.700001n V_hig
+ 37.800000n V_hig
+ 37.800001n V_hig
+ 37.900000n V_hig
+ 37.900001n V_hig
+ 38.000000n V_hig
+ 38.000001n V_low
+ 38.100000n V_low
+ 38.100001n V_low
+ 38.200000n V_low
+ 38.200001n V_low
+ 38.300000n V_low
+ 38.300001n V_low
+ 38.400000n V_low
+ 38.400001n V_low
+ 38.500000n V_low
+ 38.500001n V_low
+ 38.600000n V_low
+ 38.600001n V_low
+ 38.700000n V_low
+ 38.700001n V_low
+ 38.800000n V_low
+ 38.800001n V_low
+ 38.900000n V_low
+ 38.900001n V_low
+ 39.000000n V_low
+ 39.000001n V_low
+ 39.100000n V_low
+ 39.100001n V_low
+ 39.200000n V_low
+ 39.200001n V_low
+ 39.300000n V_low
+ 39.300001n V_low
+ 39.400000n V_low
+ 39.400001n V_low
+ 39.500000n V_low
+ 39.500001n V_low
+ 39.600000n V_low
+ 39.600001n V_low
+ 39.700000n V_low
+ 39.700001n V_low
+ 39.800000n V_low
+ 39.800001n V_low
+ 39.900000n V_low
+ 39.900001n V_low
+ 40.000000n V_low
+ 40.000001n V_hig
+ 40.100000n V_hig
+ 40.100001n V_hig
+ 40.200000n V_hig
+ 40.200001n V_hig
+ 40.300000n V_hig
+ 40.300001n V_hig
+ 40.400000n V_hig
+ 40.400001n V_hig
+ 40.500000n V_hig
+ 40.500001n V_hig
+ 40.600000n V_hig
+ 40.600001n V_hig
+ 40.700000n V_hig
+ 40.700001n V_hig
+ 40.800000n V_hig
+ 40.800001n V_hig
+ 40.900000n V_hig
+ 40.900001n V_hig
+ 41.000000n V_hig
+ 41.000001n V_hig
+ 41.100000n V_hig
+ 41.100001n V_hig
+ 41.200000n V_hig
+ 41.200001n V_hig
+ 41.300000n V_hig
+ 41.300001n V_hig
+ 41.400000n V_hig
+ 41.400001n V_hig
+ 41.500000n V_hig
+ 41.500001n V_hig
+ 41.600000n V_hig
+ 41.600001n V_hig
+ 41.700000n V_hig
+ 41.700001n V_hig
+ 41.800000n V_hig
+ 41.800001n V_hig
+ 41.900000n V_hig
+ 41.900001n V_hig
+ 42.000000n V_hig
+ 42.000001n V_hig
+ 42.100000n V_hig
+ 42.100001n V_hig
+ 42.200000n V_hig
+ 42.200001n V_hig
+ 42.300000n V_hig
+ 42.300001n V_hig
+ 42.400000n V_hig
+ 42.400001n V_hig
+ 42.500000n V_hig
+ 42.500001n V_hig
+ 42.600000n V_hig
+ 42.600001n V_hig
+ 42.700000n V_hig
+ 42.700001n V_hig
+ 42.800000n V_hig
+ 42.800001n V_hig
+ 42.900000n V_hig
+ 42.900001n V_hig
+ 43.000000n V_hig
+ 43.000001n V_low
+ 43.100000n V_low
+ 43.100001n V_low
+ 43.200000n V_low
+ 43.200001n V_low
+ 43.300000n V_low
+ 43.300001n V_low
+ 43.400000n V_low
+ 43.400001n V_low
+ 43.500000n V_low
+ 43.500001n V_low
+ 43.600000n V_low
+ 43.600001n V_low
+ 43.700000n V_low
+ 43.700001n V_low
+ 43.800000n V_low
+ 43.800001n V_low
+ 43.900000n V_low
+ 43.900001n V_low
+ 44.000000n V_low
+ 44.000001n V_hig
+ 44.100000n V_hig
+ 44.100001n V_hig
+ 44.200000n V_hig
+ 44.200001n V_hig
+ 44.300000n V_hig
+ 44.300001n V_hig
+ 44.400000n V_hig
+ 44.400001n V_hig
+ 44.500000n V_hig
+ 44.500001n V_hig
+ 44.600000n V_hig
+ 44.600001n V_hig
+ 44.700000n V_hig
+ 44.700001n V_hig
+ 44.800000n V_hig
+ 44.800001n V_hig
+ 44.900000n V_hig
+ 44.900001n V_hig
+ 45.000000n V_hig
+ 45.000001n V_hig
+ 45.100000n V_hig
+ 45.100001n V_hig
+ 45.200000n V_hig
+ 45.200001n V_hig
+ 45.300000n V_hig
+ 45.300001n V_hig
+ 45.400000n V_hig
+ 45.400001n V_hig
+ 45.500000n V_hig
+ 45.500001n V_hig
+ 45.600000n V_hig
+ 45.600001n V_hig
+ 45.700000n V_hig
+ 45.700001n V_hig
+ 45.800000n V_hig
+ 45.800001n V_hig
+ 45.900000n V_hig
+ 45.900001n V_hig
+ 46.000000n V_hig
+ 46.000001n V_low
+ 46.100000n V_low
+ 46.100001n V_low
+ 46.200000n V_low
+ 46.200001n V_low
+ 46.300000n V_low
+ 46.300001n V_low
+ 46.400000n V_low
+ 46.400001n V_low
+ 46.500000n V_low
+ 46.500001n V_low
+ 46.600000n V_low
+ 46.600001n V_low
+ 46.700000n V_low
+ 46.700001n V_low
+ 46.800000n V_low
+ 46.800001n V_low
+ 46.900000n V_low
+ 46.900001n V_low
+ 47.000000n V_low
+ 47.000001n V_hig
+ 47.100000n V_hig
+ 47.100001n V_hig
+ 47.200000n V_hig
+ 47.200001n V_hig
+ 47.300000n V_hig
+ 47.300001n V_hig
+ 47.400000n V_hig
+ 47.400001n V_hig
+ 47.500000n V_hig
+ 47.500001n V_hig
+ 47.600000n V_hig
+ 47.600001n V_hig
+ 47.700000n V_hig
+ 47.700001n V_hig
+ 47.800000n V_hig
+ 47.800001n V_hig
+ 47.900000n V_hig
+ 47.900001n V_hig
+ 48.000000n V_hig
+ 48.000001n V_hig
+ 48.100000n V_hig
+ 48.100001n V_hig
+ 48.200000n V_hig
+ 48.200001n V_hig
+ 48.300000n V_hig
+ 48.300001n V_hig
+ 48.400000n V_hig
+ 48.400001n V_hig
+ 48.500000n V_hig
+ 48.500001n V_hig
+ 48.600000n V_hig
+ 48.600001n V_hig
+ 48.700000n V_hig
+ 48.700001n V_hig
+ 48.800000n V_hig
+ 48.800001n V_hig
+ 48.900000n V_hig
+ 48.900001n V_hig
+ 49.000000n V_hig
+ 49.000001n V_low
+ 49.100000n V_low
+ 49.100001n V_low
+ 49.200000n V_low
+ 49.200001n V_low
+ 49.300000n V_low
+ 49.300001n V_low
+ 49.400000n V_low
+ 49.400001n V_low
+ 49.500000n V_low
+ 49.500001n V_low
+ 49.600000n V_low
+ 49.600001n V_low
+ 49.700000n V_low
+ 49.700001n V_low
+ 49.800000n V_low
+ 49.800001n V_low
+ 49.900000n V_low
+ 49.900001n V_low
+ 50.000000n V_low
+ 50.000001n V_low
+ 50.100000n V_low
+ 50.100001n V_low
+ 50.200000n V_low
+ 50.200001n V_low
+ 50.300000n V_low
+ 50.300001n V_low
+ 50.400000n V_low
+ 50.400001n V_low
+ 50.500000n V_low
+ 50.500001n V_low
+ 50.600000n V_low
+ 50.600001n V_low
+ 50.700000n V_low
+ 50.700001n V_low
+ 50.800000n V_low
+ 50.800001n V_low
+ 50.900000n V_low
+ 50.900001n V_low
+ 51.000000n V_low
+ 51.000001n V_low
+ 51.100000n V_low
+ 51.100001n V_low
+ 51.200000n V_low
+ 51.200001n V_low
+ 51.300000n V_low
+ 51.300001n V_low
+ 51.400000n V_low
+ 51.400001n V_low
+ 51.500000n V_low
+ 51.500001n V_low
+ 51.600000n V_low
+ 51.600001n V_low
+ 51.700000n V_low
+ 51.700001n V_low
+ 51.800000n V_low
+ 51.800001n V_low
+ 51.900000n V_low
+ 51.900001n V_low
+ 52.000000n V_low
+ 52.000001n V_hig
+ 52.100000n V_hig
+ 52.100001n V_hig
+ 52.200000n V_hig
+ 52.200001n V_hig
+ 52.300000n V_hig
+ 52.300001n V_hig
+ 52.400000n V_hig
+ 52.400001n V_hig
+ 52.500000n V_hig
+ 52.500001n V_hig
+ 52.600000n V_hig
+ 52.600001n V_hig
+ 52.700000n V_hig
+ 52.700001n V_hig
+ 52.800000n V_hig
+ 52.800001n V_hig
+ 52.900000n V_hig
+ 52.900001n V_hig
+ 53.000000n V_hig
+ 53.000001n V_hig
+ 53.100000n V_hig
+ 53.100001n V_hig
+ 53.200000n V_hig
+ 53.200001n V_hig
+ 53.300000n V_hig
+ 53.300001n V_hig
+ 53.400000n V_hig
+ 53.400001n V_hig
+ 53.500000n V_hig
+ 53.500001n V_hig
+ 53.600000n V_hig
+ 53.600001n V_hig
+ 53.700000n V_hig
+ 53.700001n V_hig
+ 53.800000n V_hig
+ 53.800001n V_hig
+ 53.900000n V_hig
+ 53.900001n V_hig
+ 54.000000n V_hig
+ 54.000001n V_low
+ 54.100000n V_low
+ 54.100001n V_low
+ 54.200000n V_low
+ 54.200001n V_low
+ 54.300000n V_low
+ 54.300001n V_low
+ 54.400000n V_low
+ 54.400001n V_low
+ 54.500000n V_low
+ 54.500001n V_low
+ 54.600000n V_low
+ 54.600001n V_low
+ 54.700000n V_low
+ 54.700001n V_low
+ 54.800000n V_low
+ 54.800001n V_low
+ 54.900000n V_low
+ 54.900001n V_low
+ 55.000000n V_low
+ 55.000001n V_low
+ 55.100000n V_low
+ 55.100001n V_low
+ 55.200000n V_low
+ 55.200001n V_low
+ 55.300000n V_low
+ 55.300001n V_low
+ 55.400000n V_low
+ 55.400001n V_low
+ 55.500000n V_low
+ 55.500001n V_low
+ 55.600000n V_low
+ 55.600001n V_low
+ 55.700000n V_low
+ 55.700001n V_low
+ 55.800000n V_low
+ 55.800001n V_low
+ 55.900000n V_low
+ 55.900001n V_low
+ 56.000000n V_low
+ 56.000001n V_hig
+ 56.100000n V_hig
+ 56.100001n V_hig
+ 56.200000n V_hig
+ 56.200001n V_hig
+ 56.300000n V_hig
+ 56.300001n V_hig
+ 56.400000n V_hig
+ 56.400001n V_hig
+ 56.500000n V_hig
+ 56.500001n V_hig
+ 56.600000n V_hig
+ 56.600001n V_hig
+ 56.700000n V_hig
+ 56.700001n V_hig
+ 56.800000n V_hig
+ 56.800001n V_hig
+ 56.900000n V_hig
+ 56.900001n V_hig
+ 57.000000n V_hig
+ 57.000001n V_low
+ 57.100000n V_low
+ 57.100001n V_low
+ 57.200000n V_low
+ 57.200001n V_low
+ 57.300000n V_low
+ 57.300001n V_low
+ 57.400000n V_low
+ 57.400001n V_low
+ 57.500000n V_low
+ 57.500001n V_low
+ 57.600000n V_low
+ 57.600001n V_low
+ 57.700000n V_low
+ 57.700001n V_low
+ 57.800000n V_low
+ 57.800001n V_low
+ 57.900000n V_low
+ 57.900001n V_low
+ 58.000000n V_low
+ 58.000001n V_hig
+ 58.100000n V_hig
+ 58.100001n V_hig
+ 58.200000n V_hig
+ 58.200001n V_hig
+ 58.300000n V_hig
+ 58.300001n V_hig
+ 58.400000n V_hig
+ 58.400001n V_hig
+ 58.500000n V_hig
+ 58.500001n V_hig
+ 58.600000n V_hig
+ 58.600001n V_hig
+ 58.700000n V_hig
+ 58.700001n V_hig
+ 58.800000n V_hig
+ 58.800001n V_hig
+ 58.900000n V_hig
+ 58.900001n V_hig
+ 59.000000n V_hig
+ 59.000001n V_low
+ 59.100000n V_low
+ 59.100001n V_low
+ 59.200000n V_low
+ 59.200001n V_low
+ 59.300000n V_low
+ 59.300001n V_low
+ 59.400000n V_low
+ 59.400001n V_low
+ 59.500000n V_low
+ 59.500001n V_low
+ 59.600000n V_low
+ 59.600001n V_low
+ 59.700000n V_low
+ 59.700001n V_low
+ 59.800000n V_low
+ 59.800001n V_low
+ 59.900000n V_low
+ 59.900001n V_low
+ 60.000000n V_low
+ 60.000001n V_low
+ 60.100000n V_low
+ 60.100001n V_low
+ 60.200000n V_low
+ 60.200001n V_low
+ 60.300000n V_low
+ 60.300001n V_low
+ 60.400000n V_low
+ 60.400001n V_low
+ 60.500000n V_low
+ 60.500001n V_low
+ 60.600000n V_low
+ 60.600001n V_low
+ 60.700000n V_low
+ 60.700001n V_low
+ 60.800000n V_low
+ 60.800001n V_low
+ 60.900000n V_low
+ 60.900001n V_low
+ 61.000000n V_low
+ 61.000001n V_low
+ 61.100000n V_low
+ 61.100001n V_low
+ 61.200000n V_low
+ 61.200001n V_low
+ 61.300000n V_low
+ 61.300001n V_low
+ 61.400000n V_low
+ 61.400001n V_low
+ 61.500000n V_low
+ 61.500001n V_low
+ 61.600000n V_low
+ 61.600001n V_low
+ 61.700000n V_low
+ 61.700001n V_low
+ 61.800000n V_low
+ 61.800001n V_low
+ 61.900000n V_low
+ 61.900001n V_low
+ 62.000000n V_low
+ 62.000001n V_hig
+ 62.100000n V_hig
+ 62.100001n V_hig
+ 62.200000n V_hig
+ 62.200001n V_hig
+ 62.300000n V_hig
+ 62.300001n V_hig
+ 62.400000n V_hig
+ 62.400001n V_hig
+ 62.500000n V_hig
+ 62.500001n V_hig
+ 62.600000n V_hig
+ 62.600001n V_hig
+ 62.700000n V_hig
+ 62.700001n V_hig
+ 62.800000n V_hig
+ 62.800001n V_hig
+ 62.900000n V_hig
+ 62.900001n V_hig
+ 63.000000n V_hig
+ 63.000001n V_low
+ 63.100000n V_low
+ 63.100001n V_low
+ 63.200000n V_low
+ 63.200001n V_low
+ 63.300000n V_low
+ 63.300001n V_low
+ 63.400000n V_low
+ 63.400001n V_low
+ 63.500000n V_low
+ 63.500001n V_low
+ 63.600000n V_low
+ 63.600001n V_low
+ 63.700000n V_low
+ 63.700001n V_low
+ 63.800000n V_low
+ 63.800001n V_low
+ 63.900000n V_low
+ 63.900001n V_low
+ 64.000000n V_low
+ 64.000001n V_low
+ 64.100000n V_low
+ 64.100001n V_low
+ 64.200000n V_low
+ 64.200001n V_low
+ 64.300000n V_low
+ 64.300001n V_low
+ 64.400000n V_low
+ 64.400001n V_low
+ 64.500000n V_low
+ 64.500001n V_low
+ 64.600000n V_low
+ 64.600001n V_low
+ 64.700000n V_low
+ 64.700001n V_low
+ 64.800000n V_low
+ 64.800001n V_low
+ 64.900000n V_low
+ 64.900001n V_low
+ 65.000000n V_low
+ 65.000001n V_low
+ 65.100000n V_low
+ 65.100001n V_low
+ 65.200000n V_low
+ 65.200001n V_low
+ 65.300000n V_low
+ 65.300001n V_low
+ 65.400000n V_low
+ 65.400001n V_low
+ 65.500000n V_low
+ 65.500001n V_low
+ 65.600000n V_low
+ 65.600001n V_low
+ 65.700000n V_low
+ 65.700001n V_low
+ 65.800000n V_low
+ 65.800001n V_low
+ 65.900000n V_low
+ 65.900001n V_low
+ 66.000000n V_low
+ 66.000001n V_hig
+ 66.100000n V_hig
+ 66.100001n V_hig
+ 66.200000n V_hig
+ 66.200001n V_hig
+ 66.300000n V_hig
+ 66.300001n V_hig
+ 66.400000n V_hig
+ 66.400001n V_hig
+ 66.500000n V_hig
+ 66.500001n V_hig
+ 66.600000n V_hig
+ 66.600001n V_hig
+ 66.700000n V_hig
+ 66.700001n V_hig
+ 66.800000n V_hig
+ 66.800001n V_hig
+ 66.900000n V_hig
+ 66.900001n V_hig
+ 67.000000n V_hig
+ 67.000001n V_low
+ 67.100000n V_low
+ 67.100001n V_low
+ 67.200000n V_low
+ 67.200001n V_low
+ 67.300000n V_low
+ 67.300001n V_low
+ 67.400000n V_low
+ 67.400001n V_low
+ 67.500000n V_low
+ 67.500001n V_low
+ 67.600000n V_low
+ 67.600001n V_low
+ 67.700000n V_low
+ 67.700001n V_low
+ 67.800000n V_low
+ 67.800001n V_low
+ 67.900000n V_low
+ 67.900001n V_low
+ 68.000000n V_low
+ 68.000001n V_hig
+ 68.100000n V_hig
+ 68.100001n V_hig
+ 68.200000n V_hig
+ 68.200001n V_hig
+ 68.300000n V_hig
+ 68.300001n V_hig
+ 68.400000n V_hig
+ 68.400001n V_hig
+ 68.500000n V_hig
+ 68.500001n V_hig
+ 68.600000n V_hig
+ 68.600001n V_hig
+ 68.700000n V_hig
+ 68.700001n V_hig
+ 68.800000n V_hig
+ 68.800001n V_hig
+ 68.900000n V_hig
+ 68.900001n V_hig
+ 69.000000n V_hig
+ 69.000001n V_low
+ 69.100000n V_low
+ 69.100001n V_low
+ 69.200000n V_low
+ 69.200001n V_low
+ 69.300000n V_low
+ 69.300001n V_low
+ 69.400000n V_low
+ 69.400001n V_low
+ 69.500000n V_low
+ 69.500001n V_low
+ 69.600000n V_low
+ 69.600001n V_low
+ 69.700000n V_low
+ 69.700001n V_low
+ 69.800000n V_low
+ 69.800001n V_low
+ 69.900000n V_low
+ 69.900001n V_low
+ 70.000000n V_low
+ 70.000001n V_hig
+ 70.100000n V_hig
+ 70.100001n V_hig
+ 70.200000n V_hig
+ 70.200001n V_hig
+ 70.300000n V_hig
+ 70.300001n V_hig
+ 70.400000n V_hig
+ 70.400001n V_hig
+ 70.500000n V_hig
+ 70.500001n V_hig
+ 70.600000n V_hig
+ 70.600001n V_hig
+ 70.700000n V_hig
+ 70.700001n V_hig
+ 70.800000n V_hig
+ 70.800001n V_hig
+ 70.900000n V_hig
+ 70.900001n V_hig
+ 71.000000n V_hig
+ 71.000001n V_hig
+ 71.100000n V_hig
+ 71.100001n V_hig
+ 71.200000n V_hig
+ 71.200001n V_hig
+ 71.300000n V_hig
+ 71.300001n V_hig
+ 71.400000n V_hig
+ 71.400001n V_hig
+ 71.500000n V_hig
+ 71.500001n V_hig
+ 71.600000n V_hig
+ 71.600001n V_hig
+ 71.700000n V_hig
+ 71.700001n V_hig
+ 71.800000n V_hig
+ 71.800001n V_hig
+ 71.900000n V_hig
+ 71.900001n V_hig
+ 72.000000n V_hig
+ 72.000001n V_low
+ 72.100000n V_low
+ 72.100001n V_low
+ 72.200000n V_low
+ 72.200001n V_low
+ 72.300000n V_low
+ 72.300001n V_low
+ 72.400000n V_low
+ 72.400001n V_low
+ 72.500000n V_low
+ 72.500001n V_low
+ 72.600000n V_low
+ 72.600001n V_low
+ 72.700000n V_low
+ 72.700001n V_low
+ 72.800000n V_low
+ 72.800001n V_low
+ 72.900000n V_low
+ 72.900001n V_low
+ 73.000000n V_low
+ 73.000001n V_low
+ 73.100000n V_low
+ 73.100001n V_low
+ 73.200000n V_low
+ 73.200001n V_low
+ 73.300000n V_low
+ 73.300001n V_low
+ 73.400000n V_low
+ 73.400001n V_low
+ 73.500000n V_low
+ 73.500001n V_low
+ 73.600000n V_low
+ 73.600001n V_low
+ 73.700000n V_low
+ 73.700001n V_low
+ 73.800000n V_low
+ 73.800001n V_low
+ 73.900000n V_low
+ 73.900001n V_low
+ 74.000000n V_low
+ 74.000001n V_hig
+ 74.100000n V_hig
+ 74.100001n V_hig
+ 74.200000n V_hig
+ 74.200001n V_hig
+ 74.300000n V_hig
+ 74.300001n V_hig
+ 74.400000n V_hig
+ 74.400001n V_hig
+ 74.500000n V_hig
+ 74.500001n V_hig
+ 74.600000n V_hig
+ 74.600001n V_hig
+ 74.700000n V_hig
+ 74.700001n V_hig
+ 74.800000n V_hig
+ 74.800001n V_hig
+ 74.900000n V_hig
+ 74.900001n V_hig
+ 75.000000n V_hig
+ 75.000001n V_low
+ 75.100000n V_low
+ 75.100001n V_low
+ 75.200000n V_low
+ 75.200001n V_low
+ 75.300000n V_low
+ 75.300001n V_low
+ 75.400000n V_low
+ 75.400001n V_low
+ 75.500000n V_low
+ 75.500001n V_low
+ 75.600000n V_low
+ 75.600001n V_low
+ 75.700000n V_low
+ 75.700001n V_low
+ 75.800000n V_low
+ 75.800001n V_low
+ 75.900000n V_low
+ 75.900001n V_low
+ 76.000000n V_low
+ 76.000001n V_low
+ 76.100000n V_low
+ 76.100001n V_low
+ 76.200000n V_low
+ 76.200001n V_low
+ 76.300000n V_low
+ 76.300001n V_low
+ 76.400000n V_low
+ 76.400001n V_low
+ 76.500000n V_low
+ 76.500001n V_low
+ 76.600000n V_low
+ 76.600001n V_low
+ 76.700000n V_low
+ 76.700001n V_low
+ 76.800000n V_low
+ 76.800001n V_low
+ 76.900000n V_low
+ 76.900001n V_low
+ 77.000000n V_low
+ 77.000001n V_low
+ 77.100000n V_low
+ 77.100001n V_low
+ 77.200000n V_low
+ 77.200001n V_low
+ 77.300000n V_low
+ 77.300001n V_low
+ 77.400000n V_low
+ 77.400001n V_low
+ 77.500000n V_low
+ 77.500001n V_low
+ 77.600000n V_low
+ 77.600001n V_low
+ 77.700000n V_low
+ 77.700001n V_low
+ 77.800000n V_low
+ 77.800001n V_low
+ 77.900000n V_low
+ 77.900001n V_low
+ 78.000000n V_low
+ 78.000001n V_low
+ 78.100000n V_low
+ 78.100001n V_low
+ 78.200000n V_low
+ 78.200001n V_low
+ 78.300000n V_low
+ 78.300001n V_low
+ 78.400000n V_low
+ 78.400001n V_low
+ 78.500000n V_low
+ 78.500001n V_low
+ 78.600000n V_low
+ 78.600001n V_low
+ 78.700000n V_low
+ 78.700001n V_low
+ 78.800000n V_low
+ 78.800001n V_low
+ 78.900000n V_low
+ 78.900001n V_low
+ 79.000000n V_low
+ 79.000001n V_hig
+ 79.100000n V_hig
+ 79.100001n V_hig
+ 79.200000n V_hig
+ 79.200001n V_hig
+ 79.300000n V_hig
+ 79.300001n V_hig
+ 79.400000n V_hig
+ 79.400001n V_hig
+ 79.500000n V_hig
+ 79.500001n V_hig
+ 79.600000n V_hig
+ 79.600001n V_hig
+ 79.700000n V_hig
+ 79.700001n V_hig
+ 79.800000n V_hig
+ 79.800001n V_hig
+ 79.900000n V_hig
+ 79.900001n V_hig
+ 80.000000n V_hig
+ 80.000001n V_hig
+ 80.100000n V_hig
+ 80.100001n V_hig
+ 80.200000n V_hig
+ 80.200001n V_hig
+ 80.300000n V_hig
+ 80.300001n V_hig
+ 80.400000n V_hig
+ 80.400001n V_hig
+ 80.500000n V_hig
+ 80.500001n V_hig
+ 80.600000n V_hig
+ 80.600001n V_hig
+ 80.700000n V_hig
+ 80.700001n V_hig
+ 80.800000n V_hig
+ 80.800001n V_hig
+ 80.900000n V_hig
+ 80.900001n V_hig
+ 81.000000n V_hig
+ 81.000001n V_hig
+ 81.100000n V_hig
+ 81.100001n V_hig
+ 81.200000n V_hig
+ 81.200001n V_hig
+ 81.300000n V_hig
+ 81.300001n V_hig
+ 81.400000n V_hig
+ 81.400001n V_hig
+ 81.500000n V_hig
+ 81.500001n V_hig
+ 81.600000n V_hig
+ 81.600001n V_hig
+ 81.700000n V_hig
+ 81.700001n V_hig
+ 81.800000n V_hig
+ 81.800001n V_hig
+ 81.900000n V_hig
+ 81.900001n V_hig
+ 82.000000n V_hig
+ 82.000001n V_low
+ 82.100000n V_low
+ 82.100001n V_low
+ 82.200000n V_low
+ 82.200001n V_low
+ 82.300000n V_low
+ 82.300001n V_low
+ 82.400000n V_low
+ 82.400001n V_low
+ 82.500000n V_low
+ 82.500001n V_low
+ 82.600000n V_low
+ 82.600001n V_low
+ 82.700000n V_low
+ 82.700001n V_low
+ 82.800000n V_low
+ 82.800001n V_low
+ 82.900000n V_low
+ 82.900001n V_low
+ 83.000000n V_low
+ 83.000001n V_low
+ 83.100000n V_low
+ 83.100001n V_low
+ 83.200000n V_low
+ 83.200001n V_low
+ 83.300000n V_low
+ 83.300001n V_low
+ 83.400000n V_low
+ 83.400001n V_low
+ 83.500000n V_low
+ 83.500001n V_low
+ 83.600000n V_low
+ 83.600001n V_low
+ 83.700000n V_low
+ 83.700001n V_low
+ 83.800000n V_low
+ 83.800001n V_low
+ 83.900000n V_low
+ 83.900001n V_low
+ 84.000000n V_low
+ 84.000001n V_low
+ 84.100000n V_low
+ 84.100001n V_low
+ 84.200000n V_low
+ 84.200001n V_low
+ 84.300000n V_low
+ 84.300001n V_low
+ 84.400000n V_low
+ 84.400001n V_low
+ 84.500000n V_low
+ 84.500001n V_low
+ 84.600000n V_low
+ 84.600001n V_low
+ 84.700000n V_low
+ 84.700001n V_low
+ 84.800000n V_low
+ 84.800001n V_low
+ 84.900000n V_low
+ 84.900001n V_low
+ 85.000000n V_low
+ 85.000001n V_hig
+ 85.100000n V_hig
+ 85.100001n V_hig
+ 85.200000n V_hig
+ 85.200001n V_hig
+ 85.300000n V_hig
+ 85.300001n V_hig
+ 85.400000n V_hig
+ 85.400001n V_hig
+ 85.500000n V_hig
+ 85.500001n V_hig
+ 85.600000n V_hig
+ 85.600001n V_hig
+ 85.700000n V_hig
+ 85.700001n V_hig
+ 85.800000n V_hig
+ 85.800001n V_hig
+ 85.900000n V_hig
+ 85.900001n V_hig
+ 86.000000n V_hig
+ 86.000001n V_hig
+ 86.100000n V_hig
+ 86.100001n V_hig
+ 86.200000n V_hig
+ 86.200001n V_hig
+ 86.300000n V_hig
+ 86.300001n V_hig
+ 86.400000n V_hig
+ 86.400001n V_hig
+ 86.500000n V_hig
+ 86.500001n V_hig
+ 86.600000n V_hig
+ 86.600001n V_hig
+ 86.700000n V_hig
+ 86.700001n V_hig
+ 86.800000n V_hig
+ 86.800001n V_hig
+ 86.900000n V_hig
+ 86.900001n V_hig
+ 87.000000n V_hig
+ 87.000001n V_low
+ 87.100000n V_low
+ 87.100001n V_low
+ 87.200000n V_low
+ 87.200001n V_low
+ 87.300000n V_low
+ 87.300001n V_low
+ 87.400000n V_low
+ 87.400001n V_low
+ 87.500000n V_low
+ 87.500001n V_low
+ 87.600000n V_low
+ 87.600001n V_low
+ 87.700000n V_low
+ 87.700001n V_low
+ 87.800000n V_low
+ 87.800001n V_low
+ 87.900000n V_low
+ 87.900001n V_low
+ 88.000000n V_low
+ 88.000001n V_hig
+ 88.100000n V_hig
+ 88.100001n V_hig
+ 88.200000n V_hig
+ 88.200001n V_hig
+ 88.300000n V_hig
+ 88.300001n V_hig
+ 88.400000n V_hig
+ 88.400001n V_hig
+ 88.500000n V_hig
+ 88.500001n V_hig
+ 88.600000n V_hig
+ 88.600001n V_hig
+ 88.700000n V_hig
+ 88.700001n V_hig
+ 88.800000n V_hig
+ 88.800001n V_hig
+ 88.900000n V_hig
+ 88.900001n V_hig
+ 89.000000n V_hig
+ 89.000001n V_low
+ 89.100000n V_low
+ 89.100001n V_low
+ 89.200000n V_low
+ 89.200001n V_low
+ 89.300000n V_low
+ 89.300001n V_low
+ 89.400000n V_low
+ 89.400001n V_low
+ 89.500000n V_low
+ 89.500001n V_low
+ 89.600000n V_low
+ 89.600001n V_low
+ 89.700000n V_low
+ 89.700001n V_low
+ 89.800000n V_low
+ 89.800001n V_low
+ 89.900000n V_low
+ 89.900001n V_low
+ 90.000000n V_low
+ 90.000001n V_hig
+ 90.100000n V_hig
+ 90.100001n V_hig
+ 90.200000n V_hig
+ 90.200001n V_hig
+ 90.300000n V_hig
+ 90.300001n V_hig
+ 90.400000n V_hig
+ 90.400001n V_hig
+ 90.500000n V_hig
+ 90.500001n V_hig
+ 90.600000n V_hig
+ 90.600001n V_hig
+ 90.700000n V_hig
+ 90.700001n V_hig
+ 90.800000n V_hig
+ 90.800001n V_hig
+ 90.900000n V_hig
+ 90.900001n V_hig
+ 91.000000n V_hig
+ 91.000001n V_hig
+ 91.100000n V_hig
+ 91.100001n V_hig
+ 91.200000n V_hig
+ 91.200001n V_hig
+ 91.300000n V_hig
+ 91.300001n V_hig
+ 91.400000n V_hig
+ 91.400001n V_hig
+ 91.500000n V_hig
+ 91.500001n V_hig
+ 91.600000n V_hig
+ 91.600001n V_hig
+ 91.700000n V_hig
+ 91.700001n V_hig
+ 91.800000n V_hig
+ 91.800001n V_hig
+ 91.900000n V_hig
+ 91.900001n V_hig
+ 92.000000n V_hig
+ 92.000001n V_low
+ 92.100000n V_low
+ 92.100001n V_low
+ 92.200000n V_low
+ 92.200001n V_low
+ 92.300000n V_low
+ 92.300001n V_low
+ 92.400000n V_low
+ 92.400001n V_low
+ 92.500000n V_low
+ 92.500001n V_low
+ 92.600000n V_low
+ 92.600001n V_low
+ 92.700000n V_low
+ 92.700001n V_low
+ 92.800000n V_low
+ 92.800001n V_low
+ 92.900000n V_low
+ 92.900001n V_low
+ 93.000000n V_low
+ 93.000001n V_hig
+ 93.100000n V_hig
+ 93.100001n V_hig
+ 93.200000n V_hig
+ 93.200001n V_hig
+ 93.300000n V_hig
+ 93.300001n V_hig
+ 93.400000n V_hig
+ 93.400001n V_hig
+ 93.500000n V_hig
+ 93.500001n V_hig
+ 93.600000n V_hig
+ 93.600001n V_hig
+ 93.700000n V_hig
+ 93.700001n V_hig
+ 93.800000n V_hig
+ 93.800001n V_hig
+ 93.900000n V_hig
+ 93.900001n V_hig
+ 94.000000n V_hig
+ 94.000001n V_low
+ 94.100000n V_low
+ 94.100001n V_low
+ 94.200000n V_low
+ 94.200001n V_low
+ 94.300000n V_low
+ 94.300001n V_low
+ 94.400000n V_low
+ 94.400001n V_low
+ 94.500000n V_low
+ 94.500001n V_low
+ 94.600000n V_low
+ 94.600001n V_low
+ 94.700000n V_low
+ 94.700001n V_low
+ 94.800000n V_low
+ 94.800001n V_low
+ 94.900000n V_low
+ 94.900001n V_low
+ 95.000000n V_low
+ 95.000001n V_hig
+ 95.100000n V_hig
+ 95.100001n V_hig
+ 95.200000n V_hig
+ 95.200001n V_hig
+ 95.300000n V_hig
+ 95.300001n V_hig
+ 95.400000n V_hig
+ 95.400001n V_hig
+ 95.500000n V_hig
+ 95.500001n V_hig
+ 95.600000n V_hig
+ 95.600001n V_hig
+ 95.700000n V_hig
+ 95.700001n V_hig
+ 95.800000n V_hig
+ 95.800001n V_hig
+ 95.900000n V_hig
+ 95.900001n V_hig
+ 96.000000n V_hig
+ 96.000001n V_hig
+ 96.100000n V_hig
+ 96.100001n V_hig
+ 96.200000n V_hig
+ 96.200001n V_hig
+ 96.300000n V_hig
+ 96.300001n V_hig
+ 96.400000n V_hig
+ 96.400001n V_hig
+ 96.500000n V_hig
+ 96.500001n V_hig
+ 96.600000n V_hig
+ 96.600001n V_hig
+ 96.700000n V_hig
+ 96.700001n V_hig
+ 96.800000n V_hig
+ 96.800001n V_hig
+ 96.900000n V_hig
+ 96.900001n V_hig
+ 97.000000n V_hig
+ 97.000001n V_low
+ 97.100000n V_low
+ 97.100001n V_low
+ 97.200000n V_low
+ 97.200001n V_low
+ 97.300000n V_low
+ 97.300001n V_low
+ 97.400000n V_low
+ 97.400001n V_low
+ 97.500000n V_low
+ 97.500001n V_low
+ 97.600000n V_low
+ 97.600001n V_low
+ 97.700000n V_low
+ 97.700001n V_low
+ 97.800000n V_low
+ 97.800001n V_low
+ 97.900000n V_low
+ 97.900001n V_low
+ 98.000000n V_low
+ 98.000001n V_hig
+ 98.100000n V_hig
+ 98.100001n V_hig
+ 98.200000n V_hig
+ 98.200001n V_hig
+ 98.300000n V_hig
+ 98.300001n V_hig
+ 98.400000n V_hig
+ 98.400001n V_hig
+ 98.500000n V_hig
+ 98.500001n V_hig
+ 98.600000n V_hig
+ 98.600001n V_hig
+ 98.700000n V_hig
+ 98.700001n V_hig
+ 98.800000n V_hig
+ 98.800001n V_hig
+ 98.900000n V_hig
+ 98.900001n V_hig
+ 99.000000n V_hig
+ 99.000001n V_low
+ 99.100000n V_low
+ 99.100001n V_low
+ 99.200000n V_low
+ 99.200001n V_low
+ 99.300000n V_low
+ 99.300001n V_low
+ 99.400000n V_low
+ 99.400001n V_low
+ 99.500000n V_low
+ 99.500001n V_low
+ 99.600000n V_low
+ 99.600001n V_low
+ 99.700000n V_low
+ 99.700001n V_low
+ 99.800000n V_low
+ 99.800001n V_low
+ 99.900000n V_low
+ 99.900001n V_low
+ 100.000000n V_low
+ 100.000001n V_low
+ 100.100000n V_low
+ 100.100001n V_low
+ 100.200000n V_low
+ 100.200001n V_low
+ 100.300000n V_low
+ 100.300001n V_low
+ 100.400000n V_low
+ 100.400001n V_low
+ 100.500000n V_low
+ 100.500001n V_low
+ 100.600000n V_low
+ 100.600001n V_low
+ 100.700000n V_low
+ 100.700001n V_low
+ 100.800000n V_low
+ 100.800001n V_low
+ 100.900000n V_low
+ 100.900001n V_low
+ 101.000000n V_low
+ 101.000001n V_hig
+ 101.100000n V_hig
+ 101.100001n V_hig
+ 101.200000n V_hig
+ 101.200001n V_hig
+ 101.300000n V_hig
+ 101.300001n V_hig
+ 101.400000n V_hig
+ 101.400001n V_hig
+ 101.500000n V_hig
+ 101.500001n V_hig
+ 101.600000n V_hig
+ 101.600001n V_hig
+ 101.700000n V_hig
+ 101.700001n V_hig
+ 101.800000n V_hig
+ 101.800001n V_hig
+ 101.900000n V_hig
+ 101.900001n V_hig
+ 102.000000n V_hig
+ 102.000001n V_low
+ 102.100000n V_low
+ 102.100001n V_low
+ 102.200000n V_low
+ 102.200001n V_low
+ 102.300000n V_low
+ 102.300001n V_low
+ 102.400000n V_low
+ 102.400001n V_low
+ 102.500000n V_low
+ 102.500001n V_low
+ 102.600000n V_low
+ 102.600001n V_low
+ 102.700000n V_low
+ 102.700001n V_low
+ 102.800000n V_low
+ 102.800001n V_low
+ 102.900000n V_low
+ 102.900001n V_low
+ 103.000000n V_low
+ 103.000001n V_hig
+ 103.100000n V_hig
+ 103.100001n V_hig
+ 103.200000n V_hig
+ 103.200001n V_hig
+ 103.300000n V_hig
+ 103.300001n V_hig
+ 103.400000n V_hig
+ 103.400001n V_hig
+ 103.500000n V_hig
+ 103.500001n V_hig
+ 103.600000n V_hig
+ 103.600001n V_hig
+ 103.700000n V_hig
+ 103.700001n V_hig
+ 103.800000n V_hig
+ 103.800001n V_hig
+ 103.900000n V_hig
+ 103.900001n V_hig
+ 104.000000n V_hig
+ 104.000001n V_hig
+ 104.100000n V_hig
+ 104.100001n V_hig
+ 104.200000n V_hig
+ 104.200001n V_hig
+ 104.300000n V_hig
+ 104.300001n V_hig
+ 104.400000n V_hig
+ 104.400001n V_hig
+ 104.500000n V_hig
+ 104.500001n V_hig
+ 104.600000n V_hig
+ 104.600001n V_hig
+ 104.700000n V_hig
+ 104.700001n V_hig
+ 104.800000n V_hig
+ 104.800001n V_hig
+ 104.900000n V_hig
+ 104.900001n V_hig
+ 105.000000n V_hig
+ 105.000001n V_low
+ 105.100000n V_low
+ 105.100001n V_low
+ 105.200000n V_low
+ 105.200001n V_low
+ 105.300000n V_low
+ 105.300001n V_low
+ 105.400000n V_low
+ 105.400001n V_low
+ 105.500000n V_low
+ 105.500001n V_low
+ 105.600000n V_low
+ 105.600001n V_low
+ 105.700000n V_low
+ 105.700001n V_low
+ 105.800000n V_low
+ 105.800001n V_low
+ 105.900000n V_low
+ 105.900001n V_low
+ 106.000000n V_low
+ 106.000001n V_low
+ 106.100000n V_low
+ 106.100001n V_low
+ 106.200000n V_low
+ 106.200001n V_low
+ 106.300000n V_low
+ 106.300001n V_low
+ 106.400000n V_low
+ 106.400001n V_low
+ 106.500000n V_low
+ 106.500001n V_low
+ 106.600000n V_low
+ 106.600001n V_low
+ 106.700000n V_low
+ 106.700001n V_low
+ 106.800000n V_low
+ 106.800001n V_low
+ 106.900000n V_low
+ 106.900001n V_low
+ 107.000000n V_low
+ 107.000001n V_hig
+ 107.100000n V_hig
+ 107.100001n V_hig
+ 107.200000n V_hig
+ 107.200001n V_hig
+ 107.300000n V_hig
+ 107.300001n V_hig
+ 107.400000n V_hig
+ 107.400001n V_hig
+ 107.500000n V_hig
+ 107.500001n V_hig
+ 107.600000n V_hig
+ 107.600001n V_hig
+ 107.700000n V_hig
+ 107.700001n V_hig
+ 107.800000n V_hig
+ 107.800001n V_hig
+ 107.900000n V_hig
+ 107.900001n V_hig
+ 108.000000n V_hig
+ 108.000001n V_hig
+ 108.100000n V_hig
+ 108.100001n V_hig
+ 108.200000n V_hig
+ 108.200001n V_hig
+ 108.300000n V_hig
+ 108.300001n V_hig
+ 108.400000n V_hig
+ 108.400001n V_hig
+ 108.500000n V_hig
+ 108.500001n V_hig
+ 108.600000n V_hig
+ 108.600001n V_hig
+ 108.700000n V_hig
+ 108.700001n V_hig
+ 108.800000n V_hig
+ 108.800001n V_hig
+ 108.900000n V_hig
+ 108.900001n V_hig
+ 109.000000n V_hig
+ 109.000001n V_hig
+ 109.100000n V_hig
+ 109.100001n V_hig
+ 109.200000n V_hig
+ 109.200001n V_hig
+ 109.300000n V_hig
+ 109.300001n V_hig
+ 109.400000n V_hig
+ 109.400001n V_hig
+ 109.500000n V_hig
+ 109.500001n V_hig
+ 109.600000n V_hig
+ 109.600001n V_hig
+ 109.700000n V_hig
+ 109.700001n V_hig
+ 109.800000n V_hig
+ 109.800001n V_hig
+ 109.900000n V_hig
+ 109.900001n V_hig
+ 110.000000n V_hig
+ 110.000001n V_hig
+ 110.100000n V_hig
+ 110.100001n V_hig
+ 110.200000n V_hig
+ 110.200001n V_hig
+ 110.300000n V_hig
+ 110.300001n V_hig
+ 110.400000n V_hig
+ 110.400001n V_hig
+ 110.500000n V_hig
+ 110.500001n V_hig
+ 110.600000n V_hig
+ 110.600001n V_hig
+ 110.700000n V_hig
+ 110.700001n V_hig
+ 110.800000n V_hig
+ 110.800001n V_hig
+ 110.900000n V_hig
+ 110.900001n V_hig
+ 111.000000n V_hig
+ 111.000001n V_hig
+ 111.100000n V_hig
+ 111.100001n V_hig
+ 111.200000n V_hig
+ 111.200001n V_hig
+ 111.300000n V_hig
+ 111.300001n V_hig
+ 111.400000n V_hig
+ 111.400001n V_hig
+ 111.500000n V_hig
+ 111.500001n V_hig
+ 111.600000n V_hig
+ 111.600001n V_hig
+ 111.700000n V_hig
+ 111.700001n V_hig
+ 111.800000n V_hig
+ 111.800001n V_hig
+ 111.900000n V_hig
+ 111.900001n V_hig
+ 112.000000n V_hig
+ 112.000001n V_hig
+ 112.100000n V_hig
+ 112.100001n V_hig
+ 112.200000n V_hig
+ 112.200001n V_hig
+ 112.300000n V_hig
+ 112.300001n V_hig
+ 112.400000n V_hig
+ 112.400001n V_hig
+ 112.500000n V_hig
+ 112.500001n V_hig
+ 112.600000n V_hig
+ 112.600001n V_hig
+ 112.700000n V_hig
+ 112.700001n V_hig
+ 112.800000n V_hig
+ 112.800001n V_hig
+ 112.900000n V_hig
+ 112.900001n V_hig
+ 113.000000n V_hig
+ 113.000001n V_low
+ 113.100000n V_low
+ 113.100001n V_low
+ 113.200000n V_low
+ 113.200001n V_low
+ 113.300000n V_low
+ 113.300001n V_low
+ 113.400000n V_low
+ 113.400001n V_low
+ 113.500000n V_low
+ 113.500001n V_low
+ 113.600000n V_low
+ 113.600001n V_low
+ 113.700000n V_low
+ 113.700001n V_low
+ 113.800000n V_low
+ 113.800001n V_low
+ 113.900000n V_low
+ 113.900001n V_low
+ 114.000000n V_low
+ 114.000001n V_hig
+ 114.100000n V_hig
+ 114.100001n V_hig
+ 114.200000n V_hig
+ 114.200001n V_hig
+ 114.300000n V_hig
+ 114.300001n V_hig
+ 114.400000n V_hig
+ 114.400001n V_hig
+ 114.500000n V_hig
+ 114.500001n V_hig
+ 114.600000n V_hig
+ 114.600001n V_hig
+ 114.700000n V_hig
+ 114.700001n V_hig
+ 114.800000n V_hig
+ 114.800001n V_hig
+ 114.900000n V_hig
+ 114.900001n V_hig
+ 115.000000n V_hig
+ 115.000001n V_low
+ 115.100000n V_low
+ 115.100001n V_low
+ 115.200000n V_low
+ 115.200001n V_low
+ 115.300000n V_low
+ 115.300001n V_low
+ 115.400000n V_low
+ 115.400001n V_low
+ 115.500000n V_low
+ 115.500001n V_low
+ 115.600000n V_low
+ 115.600001n V_low
+ 115.700000n V_low
+ 115.700001n V_low
+ 115.800000n V_low
+ 115.800001n V_low
+ 115.900000n V_low
+ 115.900001n V_low
+ 116.000000n V_low
+ 116.000001n V_hig
+ 116.100000n V_hig
+ 116.100001n V_hig
+ 116.200000n V_hig
+ 116.200001n V_hig
+ 116.300000n V_hig
+ 116.300001n V_hig
+ 116.400000n V_hig
+ 116.400001n V_hig
+ 116.500000n V_hig
+ 116.500001n V_hig
+ 116.600000n V_hig
+ 116.600001n V_hig
+ 116.700000n V_hig
+ 116.700001n V_hig
+ 116.800000n V_hig
+ 116.800001n V_hig
+ 116.900000n V_hig
+ 116.900001n V_hig
+ 117.000000n V_hig
+ 117.000001n V_hig
+ 117.100000n V_hig
+ 117.100001n V_hig
+ 117.200000n V_hig
+ 117.200001n V_hig
+ 117.300000n V_hig
+ 117.300001n V_hig
+ 117.400000n V_hig
+ 117.400001n V_hig
+ 117.500000n V_hig
+ 117.500001n V_hig
+ 117.600000n V_hig
+ 117.600001n V_hig
+ 117.700000n V_hig
+ 117.700001n V_hig
+ 117.800000n V_hig
+ 117.800001n V_hig
+ 117.900000n V_hig
+ 117.900001n V_hig
+ 118.000000n V_hig
+ 118.000001n V_hig
+ 118.100000n V_hig
+ 118.100001n V_hig
+ 118.200000n V_hig
+ 118.200001n V_hig
+ 118.300000n V_hig
+ 118.300001n V_hig
+ 118.400000n V_hig
+ 118.400001n V_hig
+ 118.500000n V_hig
+ 118.500001n V_hig
+ 118.600000n V_hig
+ 118.600001n V_hig
+ 118.700000n V_hig
+ 118.700001n V_hig
+ 118.800000n V_hig
+ 118.800001n V_hig
+ 118.900000n V_hig
+ 118.900001n V_hig
+ 119.000000n V_hig
+ 119.000001n V_low
+ 119.100000n V_low
+ 119.100001n V_low
+ 119.200000n V_low
+ 119.200001n V_low
+ 119.300000n V_low
+ 119.300001n V_low
+ 119.400000n V_low
+ 119.400001n V_low
+ 119.500000n V_low
+ 119.500001n V_low
+ 119.600000n V_low
+ 119.600001n V_low
+ 119.700000n V_low
+ 119.700001n V_low
+ 119.800000n V_low
+ 119.800001n V_low
+ 119.900000n V_low
+ 119.900001n V_low
+ 120.000000n V_low
+ 120.000001n V_low
+ 120.100000n V_low
+ 120.100001n V_low
+ 120.200000n V_low
+ 120.200001n V_low
+ 120.300000n V_low
+ 120.300001n V_low
+ 120.400000n V_low
+ 120.400001n V_low
+ 120.500000n V_low
+ 120.500001n V_low
+ 120.600000n V_low
+ 120.600001n V_low
+ 120.700000n V_low
+ 120.700001n V_low
+ 120.800000n V_low
+ 120.800001n V_low
+ 120.900000n V_low
+ 120.900001n V_low
+ 121.000000n V_low
+ 121.000001n V_low
+ 121.100000n V_low
+ 121.100001n V_low
+ 121.200000n V_low
+ 121.200001n V_low
+ 121.300000n V_low
+ 121.300001n V_low
+ 121.400000n V_low
+ 121.400001n V_low
+ 121.500000n V_low
+ 121.500001n V_low
+ 121.600000n V_low
+ 121.600001n V_low
+ 121.700000n V_low
+ 121.700001n V_low
+ 121.800000n V_low
+ 121.800001n V_low
+ 121.900000n V_low
+ 121.900001n V_low
+ 122.000000n V_low
+ 122.000001n V_hig
+ 122.100000n V_hig
+ 122.100001n V_hig
+ 122.200000n V_hig
+ 122.200001n V_hig
+ 122.300000n V_hig
+ 122.300001n V_hig
+ 122.400000n V_hig
+ 122.400001n V_hig
+ 122.500000n V_hig
+ 122.500001n V_hig
+ 122.600000n V_hig
+ 122.600001n V_hig
+ 122.700000n V_hig
+ 122.700001n V_hig
+ 122.800000n V_hig
+ 122.800001n V_hig
+ 122.900000n V_hig
+ 122.900001n V_hig
+ 123.000000n V_hig
+ 123.000001n V_hig
+ 123.100000n V_hig
+ 123.100001n V_hig
+ 123.200000n V_hig
+ 123.200001n V_hig
+ 123.300000n V_hig
+ 123.300001n V_hig
+ 123.400000n V_hig
+ 123.400001n V_hig
+ 123.500000n V_hig
+ 123.500001n V_hig
+ 123.600000n V_hig
+ 123.600001n V_hig
+ 123.700000n V_hig
+ 123.700001n V_hig
+ 123.800000n V_hig
+ 123.800001n V_hig
+ 123.900000n V_hig
+ 123.900001n V_hig
+ 124.000000n V_hig
+ 124.000001n V_hig
+ 124.100000n V_hig
+ 124.100001n V_hig
+ 124.200000n V_hig
+ 124.200001n V_hig
+ 124.300000n V_hig
+ 124.300001n V_hig
+ 124.400000n V_hig
+ 124.400001n V_hig
+ 124.500000n V_hig
+ 124.500001n V_hig
+ 124.600000n V_hig
+ 124.600001n V_hig
+ 124.700000n V_hig
+ 124.700001n V_hig
+ 124.800000n V_hig
+ 124.800001n V_hig
+ 124.900000n V_hig
+ 124.900001n V_hig
+ 125.000000n V_hig
+ 125.000001n V_hig
+ 125.100000n V_hig
+ 125.100001n V_hig
+ 125.200000n V_hig
+ 125.200001n V_hig
+ 125.300000n V_hig
+ 125.300001n V_hig
+ 125.400000n V_hig
+ 125.400001n V_hig
+ 125.500000n V_hig
+ 125.500001n V_hig
+ 125.600000n V_hig
+ 125.600001n V_hig
+ 125.700000n V_hig
+ 125.700001n V_hig
+ 125.800000n V_hig
+ 125.800001n V_hig
+ 125.900000n V_hig
+ 125.900001n V_hig
+ 126.000000n V_hig
+ 126.000001n V_low
+ 126.100000n V_low
+ 126.100001n V_low
+ 126.200000n V_low
+ 126.200001n V_low
+ 126.300000n V_low
+ 126.300001n V_low
+ 126.400000n V_low
+ 126.400001n V_low
+ 126.500000n V_low
+ 126.500001n V_low
+ 126.600000n V_low
+ 126.600001n V_low
+ 126.700000n V_low
+ 126.700001n V_low
+ 126.800000n V_low
+ 126.800001n V_low
+ 126.900000n V_low
+ 126.900001n V_low
+ 127.000000n V_low
+ 127.000001n V_hig
+ 127.100000n V_hig
+ 127.100001n V_hig
+ 127.200000n V_hig
+ 127.200001n V_hig
+ 127.300000n V_hig
+ 127.300001n V_hig
+ 127.400000n V_hig
+ 127.400001n V_hig
+ 127.500000n V_hig
+ 127.500001n V_hig
+ 127.600000n V_hig
+ 127.600001n V_hig
+ 127.700000n V_hig
+ 127.700001n V_hig
+ 127.800000n V_hig
+ 127.800001n V_hig
+ 127.900000n V_hig
+ 127.900001n V_hig
+ 128.000000n V_hig
+ 128.000001n V_hig
+ 128.100000n V_hig
+ 128.100001n V_hig
+ 128.200000n V_hig
+ 128.200001n V_hig
+ 128.300000n V_hig
+ 128.300001n V_hig
+ 128.400000n V_hig
+ 128.400001n V_hig
+ 128.500000n V_hig
+ 128.500001n V_hig
+ 128.600000n V_hig
+ 128.600001n V_hig
+ 128.700000n V_hig
+ 128.700001n V_hig
+ 128.800000n V_hig
+ 128.800001n V_hig
+ 128.900000n V_hig
+ 128.900001n V_hig
+ 129.000000n V_hig
+ 129.000001n V_low
+ 129.100000n V_low
+ 129.100001n V_low
+ 129.200000n V_low
+ 129.200001n V_low
+ 129.300000n V_low
+ 129.300001n V_low
+ 129.400000n V_low
+ 129.400001n V_low
+ 129.500000n V_low
+ 129.500001n V_low
+ 129.600000n V_low
+ 129.600001n V_low
+ 129.700000n V_low
+ 129.700001n V_low
+ 129.800000n V_low
+ 129.800001n V_low
+ 129.900000n V_low
+ 129.900001n V_low
+ 130.000000n V_low
+ 130.000001n V_hig
+ 130.100000n V_hig
+ 130.100001n V_hig
+ 130.200000n V_hig
+ 130.200001n V_hig
+ 130.300000n V_hig
+ 130.300001n V_hig
+ 130.400000n V_hig
+ 130.400001n V_hig
+ 130.500000n V_hig
+ 130.500001n V_hig
+ 130.600000n V_hig
+ 130.600001n V_hig
+ 130.700000n V_hig
+ 130.700001n V_hig
+ 130.800000n V_hig
+ 130.800001n V_hig
+ 130.900000n V_hig
+ 130.900001n V_hig
+ 131.000000n V_hig
+ 131.000001n V_hig
+ 131.100000n V_hig
+ 131.100001n V_hig
+ 131.200000n V_hig
+ 131.200001n V_hig
+ 131.300000n V_hig
+ 131.300001n V_hig
+ 131.400000n V_hig
+ 131.400001n V_hig
+ 131.500000n V_hig
+ 131.500001n V_hig
+ 131.600000n V_hig
+ 131.600001n V_hig
+ 131.700000n V_hig
+ 131.700001n V_hig
+ 131.800000n V_hig
+ 131.800001n V_hig
+ 131.900000n V_hig
+ 131.900001n V_hig
+ 132.000000n V_hig
+ 132.000001n V_low
+ 132.100000n V_low
+ 132.100001n V_low
+ 132.200000n V_low
+ 132.200001n V_low
+ 132.300000n V_low
+ 132.300001n V_low
+ 132.400000n V_low
+ 132.400001n V_low
+ 132.500000n V_low
+ 132.500001n V_low
+ 132.600000n V_low
+ 132.600001n V_low
+ 132.700000n V_low
+ 132.700001n V_low
+ 132.800000n V_low
+ 132.800001n V_low
+ 132.900000n V_low
+ 132.900001n V_low
+ 133.000000n V_low
+ 133.000001n V_low
+ 133.100000n V_low
+ 133.100001n V_low
+ 133.200000n V_low
+ 133.200001n V_low
+ 133.300000n V_low
+ 133.300001n V_low
+ 133.400000n V_low
+ 133.400001n V_low
+ 133.500000n V_low
+ 133.500001n V_low
+ 133.600000n V_low
+ 133.600001n V_low
+ 133.700000n V_low
+ 133.700001n V_low
+ 133.800000n V_low
+ 133.800001n V_low
+ 133.900000n V_low
+ 133.900001n V_low
+ 134.000000n V_low
+ 134.000001n V_hig
+ 134.100000n V_hig
+ 134.100001n V_hig
+ 134.200000n V_hig
+ 134.200001n V_hig
+ 134.300000n V_hig
+ 134.300001n V_hig
+ 134.400000n V_hig
+ 134.400001n V_hig
+ 134.500000n V_hig
+ 134.500001n V_hig
+ 134.600000n V_hig
+ 134.600001n V_hig
+ 134.700000n V_hig
+ 134.700001n V_hig
+ 134.800000n V_hig
+ 134.800001n V_hig
+ 134.900000n V_hig
+ 134.900001n V_hig
+ 135.000000n V_hig
+ 135.000001n V_low
+ 135.100000n V_low
+ 135.100001n V_low
+ 135.200000n V_low
+ 135.200001n V_low
+ 135.300000n V_low
+ 135.300001n V_low
+ 135.400000n V_low
+ 135.400001n V_low
+ 135.500000n V_low
+ 135.500001n V_low
+ 135.600000n V_low
+ 135.600001n V_low
+ 135.700000n V_low
+ 135.700001n V_low
+ 135.800000n V_low
+ 135.800001n V_low
+ 135.900000n V_low
+ 135.900001n V_low
+ 136.000000n V_low
+ 136.000001n V_hig
+ 136.100000n V_hig
+ 136.100001n V_hig
+ 136.200000n V_hig
+ 136.200001n V_hig
+ 136.300000n V_hig
+ 136.300001n V_hig
+ 136.400000n V_hig
+ 136.400001n V_hig
+ 136.500000n V_hig
+ 136.500001n V_hig
+ 136.600000n V_hig
+ 136.600001n V_hig
+ 136.700000n V_hig
+ 136.700001n V_hig
+ 136.800000n V_hig
+ 136.800001n V_hig
+ 136.900000n V_hig
+ 136.900001n V_hig
+ 137.000000n V_hig
+ 137.000001n V_hig
+ 137.100000n V_hig
+ 137.100001n V_hig
+ 137.200000n V_hig
+ 137.200001n V_hig
+ 137.300000n V_hig
+ 137.300001n V_hig
+ 137.400000n V_hig
+ 137.400001n V_hig
+ 137.500000n V_hig
+ 137.500001n V_hig
+ 137.600000n V_hig
+ 137.600001n V_hig
+ 137.700000n V_hig
+ 137.700001n V_hig
+ 137.800000n V_hig
+ 137.800001n V_hig
+ 137.900000n V_hig
+ 137.900001n V_hig
+ 138.000000n V_hig
+ 138.000001n V_low
+ 138.100000n V_low
+ 138.100001n V_low
+ 138.200000n V_low
+ 138.200001n V_low
+ 138.300000n V_low
+ 138.300001n V_low
+ 138.400000n V_low
+ 138.400001n V_low
+ 138.500000n V_low
+ 138.500001n V_low
+ 138.600000n V_low
+ 138.600001n V_low
+ 138.700000n V_low
+ 138.700001n V_low
+ 138.800000n V_low
+ 138.800001n V_low
+ 138.900000n V_low
+ 138.900001n V_low
+ 139.000000n V_low
+ 139.000001n V_hig
+ 139.100000n V_hig
+ 139.100001n V_hig
+ 139.200000n V_hig
+ 139.200001n V_hig
+ 139.300000n V_hig
+ 139.300001n V_hig
+ 139.400000n V_hig
+ 139.400001n V_hig
+ 139.500000n V_hig
+ 139.500001n V_hig
+ 139.600000n V_hig
+ 139.600001n V_hig
+ 139.700000n V_hig
+ 139.700001n V_hig
+ 139.800000n V_hig
+ 139.800001n V_hig
+ 139.900000n V_hig
+ 139.900001n V_hig
+ 140.000000n V_hig
+ 140.000001n V_low
+ 140.100000n V_low
+ 140.100001n V_low
+ 140.200000n V_low
+ 140.200001n V_low
+ 140.300000n V_low
+ 140.300001n V_low
+ 140.400000n V_low
+ 140.400001n V_low
+ 140.500000n V_low
+ 140.500001n V_low
+ 140.600000n V_low
+ 140.600001n V_low
+ 140.700000n V_low
+ 140.700001n V_low
+ 140.800000n V_low
+ 140.800001n V_low
+ 140.900000n V_low
+ 140.900001n V_low
+ 141.000000n V_low
+ 141.000001n V_hig
+ 141.100000n V_hig
+ 141.100001n V_hig
+ 141.200000n V_hig
+ 141.200001n V_hig
+ 141.300000n V_hig
+ 141.300001n V_hig
+ 141.400000n V_hig
+ 141.400001n V_hig
+ 141.500000n V_hig
+ 141.500001n V_hig
+ 141.600000n V_hig
+ 141.600001n V_hig
+ 141.700000n V_hig
+ 141.700001n V_hig
+ 141.800000n V_hig
+ 141.800001n V_hig
+ 141.900000n V_hig
+ 141.900001n V_hig
+ 142.000000n V_hig
+ 142.000001n V_low
+ 142.100000n V_low
+ 142.100001n V_low
+ 142.200000n V_low
+ 142.200001n V_low
+ 142.300000n V_low
+ 142.300001n V_low
+ 142.400000n V_low
+ 142.400001n V_low
+ 142.500000n V_low
+ 142.500001n V_low
+ 142.600000n V_low
+ 142.600001n V_low
+ 142.700000n V_low
+ 142.700001n V_low
+ 142.800000n V_low
+ 142.800001n V_low
+ 142.900000n V_low
+ 142.900001n V_low
+ 143.000000n V_low
+ 143.000001n V_low
+ 143.100000n V_low
+ 143.100001n V_low
+ 143.200000n V_low
+ 143.200001n V_low
+ 143.300000n V_low
+ 143.300001n V_low
+ 143.400000n V_low
+ 143.400001n V_low
+ 143.500000n V_low
+ 143.500001n V_low
+ 143.600000n V_low
+ 143.600001n V_low
+ 143.700000n V_low
+ 143.700001n V_low
+ 143.800000n V_low
+ 143.800001n V_low
+ 143.900000n V_low
+ 143.900001n V_low
+ 144.000000n V_low
+ 144.000001n V_low
+ 144.100000n V_low
+ 144.100001n V_low
+ 144.200000n V_low
+ 144.200001n V_low
+ 144.300000n V_low
+ 144.300001n V_low
+ 144.400000n V_low
+ 144.400001n V_low
+ 144.500000n V_low
+ 144.500001n V_low
+ 144.600000n V_low
+ 144.600001n V_low
+ 144.700000n V_low
+ 144.700001n V_low
+ 144.800000n V_low
+ 144.800001n V_low
+ 144.900000n V_low
+ 144.900001n V_low
+ 145.000000n V_low
+ 145.000001n V_low
+ 145.100000n V_low
+ 145.100001n V_low
+ 145.200000n V_low
+ 145.200001n V_low
+ 145.300000n V_low
+ 145.300001n V_low
+ 145.400000n V_low
+ 145.400001n V_low
+ 145.500000n V_low
+ 145.500001n V_low
+ 145.600000n V_low
+ 145.600001n V_low
+ 145.700000n V_low
+ 145.700001n V_low
+ 145.800000n V_low
+ 145.800001n V_low
+ 145.900000n V_low
+ 145.900001n V_low
+ 146.000000n V_low
+ 146.000001n V_hig
+ 146.100000n V_hig
+ 146.100001n V_hig
+ 146.200000n V_hig
+ 146.200001n V_hig
+ 146.300000n V_hig
+ 146.300001n V_hig
+ 146.400000n V_hig
+ 146.400001n V_hig
+ 146.500000n V_hig
+ 146.500001n V_hig
+ 146.600000n V_hig
+ 146.600001n V_hig
+ 146.700000n V_hig
+ 146.700001n V_hig
+ 146.800000n V_hig
+ 146.800001n V_hig
+ 146.900000n V_hig
+ 146.900001n V_hig
+ 147.000000n V_hig
+ 147.000001n V_low
+ 147.100000n V_low
+ 147.100001n V_low
+ 147.200000n V_low
+ 147.200001n V_low
+ 147.300000n V_low
+ 147.300001n V_low
+ 147.400000n V_low
+ 147.400001n V_low
+ 147.500000n V_low
+ 147.500001n V_low
+ 147.600000n V_low
+ 147.600001n V_low
+ 147.700000n V_low
+ 147.700001n V_low
+ 147.800000n V_low
+ 147.800001n V_low
+ 147.900000n V_low
+ 147.900001n V_low
+ 148.000000n V_low
+ 148.000001n V_low
+ 148.100000n V_low
+ 148.100001n V_low
+ 148.200000n V_low
+ 148.200001n V_low
+ 148.300000n V_low
+ 148.300001n V_low
+ 148.400000n V_low
+ 148.400001n V_low
+ 148.500000n V_low
+ 148.500001n V_low
+ 148.600000n V_low
+ 148.600001n V_low
+ 148.700000n V_low
+ 148.700001n V_low
+ 148.800000n V_low
+ 148.800001n V_low
+ 148.900000n V_low
+ 148.900001n V_low
+ 149.000000n V_low
+ 149.000001n V_hig
+ 149.100000n V_hig
+ 149.100001n V_hig
+ 149.200000n V_hig
+ 149.200001n V_hig
+ 149.300000n V_hig
+ 149.300001n V_hig
+ 149.400000n V_hig
+ 149.400001n V_hig
+ 149.500000n V_hig
+ 149.500001n V_hig
+ 149.600000n V_hig
+ 149.600001n V_hig
+ 149.700000n V_hig
+ 149.700001n V_hig
+ 149.800000n V_hig
+ 149.800001n V_hig
+ 149.900000n V_hig
+ 149.900001n V_hig
+ 150.000000n V_hig
+ 150.000001n V_hig
+ 150.100000n V_hig
+ 150.100001n V_hig
+ 150.200000n V_hig
+ 150.200001n V_hig
+ 150.300000n V_hig
+ 150.300001n V_hig
+ 150.400000n V_hig
+ 150.400001n V_hig
+ 150.500000n V_hig
+ 150.500001n V_hig
+ 150.600000n V_hig
+ 150.600001n V_hig
+ 150.700000n V_hig
+ 150.700001n V_hig
+ 150.800000n V_hig
+ 150.800001n V_hig
+ 150.900000n V_hig
+ 150.900001n V_hig
+ 151.000000n V_hig
+ 151.000001n V_low
+ 151.100000n V_low
+ 151.100001n V_low
+ 151.200000n V_low
+ 151.200001n V_low
+ 151.300000n V_low
+ 151.300001n V_low
+ 151.400000n V_low
+ 151.400001n V_low
+ 151.500000n V_low
+ 151.500001n V_low
+ 151.600000n V_low
+ 151.600001n V_low
+ 151.700000n V_low
+ 151.700001n V_low
+ 151.800000n V_low
+ 151.800001n V_low
+ 151.900000n V_low
+ 151.900001n V_low
+ 152.000000n V_low
+ 152.000001n V_low
+ 152.100000n V_low
+ 152.100001n V_low
+ 152.200000n V_low
+ 152.200001n V_low
+ 152.300000n V_low
+ 152.300001n V_low
+ 152.400000n V_low
+ 152.400001n V_low
+ 152.500000n V_low
+ 152.500001n V_low
+ 152.600000n V_low
+ 152.600001n V_low
+ 152.700000n V_low
+ 152.700001n V_low
+ 152.800000n V_low
+ 152.800001n V_low
+ 152.900000n V_low
+ 152.900001n V_low
+ 153.000000n V_low
+ 153.000001n V_low
+ 153.100000n V_low
+ 153.100001n V_low
+ 153.200000n V_low
+ 153.200001n V_low
+ 153.300000n V_low
+ 153.300001n V_low
+ 153.400000n V_low
+ 153.400001n V_low
+ 153.500000n V_low
+ 153.500001n V_low
+ 153.600000n V_low
+ 153.600001n V_low
+ 153.700000n V_low
+ 153.700001n V_low
+ 153.800000n V_low
+ 153.800001n V_low
+ 153.900000n V_low
+ 153.900001n V_low
+ 154.000000n V_low
+ 154.000001n V_low
+ 154.100000n V_low
+ 154.100001n V_low
+ 154.200000n V_low
+ 154.200001n V_low
+ 154.300000n V_low
+ 154.300001n V_low
+ 154.400000n V_low
+ 154.400001n V_low
+ 154.500000n V_low
+ 154.500001n V_low
+ 154.600000n V_low
+ 154.600001n V_low
+ 154.700000n V_low
+ 154.700001n V_low
+ 154.800000n V_low
+ 154.800001n V_low
+ 154.900000n V_low
+ 154.900001n V_low
+ 155.000000n V_low
+ 155.000001n V_low
+ 155.100000n V_low
+ 155.100001n V_low
+ 155.200000n V_low
+ 155.200001n V_low
+ 155.300000n V_low
+ 155.300001n V_low
+ 155.400000n V_low
+ 155.400001n V_low
+ 155.500000n V_low
+ 155.500001n V_low
+ 155.600000n V_low
+ 155.600001n V_low
+ 155.700000n V_low
+ 155.700001n V_low
+ 155.800000n V_low
+ 155.800001n V_low
+ 155.900000n V_low
+ 155.900001n V_low
+ 156.000000n V_low
+ 156.000001n V_low
+ 156.100000n V_low
+ 156.100001n V_low
+ 156.200000n V_low
+ 156.200001n V_low
+ 156.300000n V_low
+ 156.300001n V_low
+ 156.400000n V_low
+ 156.400001n V_low
+ 156.500000n V_low
+ 156.500001n V_low
+ 156.600000n V_low
+ 156.600001n V_low
+ 156.700000n V_low
+ 156.700001n V_low
+ 156.800000n V_low
+ 156.800001n V_low
+ 156.900000n V_low
+ 156.900001n V_low
+ 157.000000n V_low
+ 157.000001n V_hig
+ 157.100000n V_hig
+ 157.100001n V_hig
+ 157.200000n V_hig
+ 157.200001n V_hig
+ 157.300000n V_hig
+ 157.300001n V_hig
+ 157.400000n V_hig
+ 157.400001n V_hig
+ 157.500000n V_hig
+ 157.500001n V_hig
+ 157.600000n V_hig
+ 157.600001n V_hig
+ 157.700000n V_hig
+ 157.700001n V_hig
+ 157.800000n V_hig
+ 157.800001n V_hig
+ 157.900000n V_hig
+ 157.900001n V_hig
+ 158.000000n V_hig
+ 158.000001n V_low
+ 158.100000n V_low
+ 158.100001n V_low
+ 158.200000n V_low
+ 158.200001n V_low
+ 158.300000n V_low
+ 158.300001n V_low
+ 158.400000n V_low
+ 158.400001n V_low
+ 158.500000n V_low
+ 158.500001n V_low
+ 158.600000n V_low
+ 158.600001n V_low
+ 158.700000n V_low
+ 158.700001n V_low
+ 158.800000n V_low
+ 158.800001n V_low
+ 158.900000n V_low
+ 158.900001n V_low
+ 159.000000n V_low
+ 159.000001n V_hig
+ 159.100000n V_hig
+ 159.100001n V_hig
+ 159.200000n V_hig
+ 159.200001n V_hig
+ 159.300000n V_hig
+ 159.300001n V_hig
+ 159.400000n V_hig
+ 159.400001n V_hig
+ 159.500000n V_hig
+ 159.500001n V_hig
+ 159.600000n V_hig
+ 159.600001n V_hig
+ 159.700000n V_hig
+ 159.700001n V_hig
+ 159.800000n V_hig
+ 159.800001n V_hig
+ 159.900000n V_hig
+ 159.900001n V_hig
+ 160.000000n V_hig
+ 160.000001n V_low
+ 160.100000n V_low
+ 160.100001n V_low
+ 160.200000n V_low
+ 160.200001n V_low
+ 160.300000n V_low
+ 160.300001n V_low
+ 160.400000n V_low
+ 160.400001n V_low
+ 160.500000n V_low
+ 160.500001n V_low
+ 160.600000n V_low
+ 160.600001n V_low
+ 160.700000n V_low
+ 160.700001n V_low
+ 160.800000n V_low
+ 160.800001n V_low
+ 160.900000n V_low
+ 160.900001n V_low
+ 161.000000n V_low
+ 161.000001n V_low
+ 161.100000n V_low
+ 161.100001n V_low
+ 161.200000n V_low
+ 161.200001n V_low
+ 161.300000n V_low
+ 161.300001n V_low
+ 161.400000n V_low
+ 161.400001n V_low
+ 161.500000n V_low
+ 161.500001n V_low
+ 161.600000n V_low
+ 161.600001n V_low
+ 161.700000n V_low
+ 161.700001n V_low
+ 161.800000n V_low
+ 161.800001n V_low
+ 161.900000n V_low
+ 161.900001n V_low
+ 162.000000n V_low
+ 162.000001n V_low
+ 162.100000n V_low
+ 162.100001n V_low
+ 162.200000n V_low
+ 162.200001n V_low
+ 162.300000n V_low
+ 162.300001n V_low
+ 162.400000n V_low
+ 162.400001n V_low
+ 162.500000n V_low
+ 162.500001n V_low
+ 162.600000n V_low
+ 162.600001n V_low
+ 162.700000n V_low
+ 162.700001n V_low
+ 162.800000n V_low
+ 162.800001n V_low
+ 162.900000n V_low
+ 162.900001n V_low
+ 163.000000n V_low
+ 163.000001n V_hig
+ 163.100000n V_hig
+ 163.100001n V_hig
+ 163.200000n V_hig
+ 163.200001n V_hig
+ 163.300000n V_hig
+ 163.300001n V_hig
+ 163.400000n V_hig
+ 163.400001n V_hig
+ 163.500000n V_hig
+ 163.500001n V_hig
+ 163.600000n V_hig
+ 163.600001n V_hig
+ 163.700000n V_hig
+ 163.700001n V_hig
+ 163.800000n V_hig
+ 163.800001n V_hig
+ 163.900000n V_hig
+ 163.900001n V_hig
+ 164.000000n V_hig
+ 164.000001n V_low
+ 164.100000n V_low
+ 164.100001n V_low
+ 164.200000n V_low
+ 164.200001n V_low
+ 164.300000n V_low
+ 164.300001n V_low
+ 164.400000n V_low
+ 164.400001n V_low
+ 164.500000n V_low
+ 164.500001n V_low
+ 164.600000n V_low
+ 164.600001n V_low
+ 164.700000n V_low
+ 164.700001n V_low
+ 164.800000n V_low
+ 164.800001n V_low
+ 164.900000n V_low
+ 164.900001n V_low
+ 165.000000n V_low
+ 165.000001n V_hig
+ 165.100000n V_hig
+ 165.100001n V_hig
+ 165.200000n V_hig
+ 165.200001n V_hig
+ 165.300000n V_hig
+ 165.300001n V_hig
+ 165.400000n V_hig
+ 165.400001n V_hig
+ 165.500000n V_hig
+ 165.500001n V_hig
+ 165.600000n V_hig
+ 165.600001n V_hig
+ 165.700000n V_hig
+ 165.700001n V_hig
+ 165.800000n V_hig
+ 165.800001n V_hig
+ 165.900000n V_hig
+ 165.900001n V_hig
+ 166.000000n V_hig
+ 166.000001n V_hig
+ 166.100000n V_hig
+ 166.100001n V_hig
+ 166.200000n V_hig
+ 166.200001n V_hig
+ 166.300000n V_hig
+ 166.300001n V_hig
+ 166.400000n V_hig
+ 166.400001n V_hig
+ 166.500000n V_hig
+ 166.500001n V_hig
+ 166.600000n V_hig
+ 166.600001n V_hig
+ 166.700000n V_hig
+ 166.700001n V_hig
+ 166.800000n V_hig
+ 166.800001n V_hig
+ 166.900000n V_hig
+ 166.900001n V_hig
+ 167.000000n V_hig
+ 167.000001n V_hig
+ 167.100000n V_hig
+ 167.100001n V_hig
+ 167.200000n V_hig
+ 167.200001n V_hig
+ 167.300000n V_hig
+ 167.300001n V_hig
+ 167.400000n V_hig
+ 167.400001n V_hig
+ 167.500000n V_hig
+ 167.500001n V_hig
+ 167.600000n V_hig
+ 167.600001n V_hig
+ 167.700000n V_hig
+ 167.700001n V_hig
+ 167.800000n V_hig
+ 167.800001n V_hig
+ 167.900000n V_hig
+ 167.900001n V_hig
+ 168.000000n V_hig
+ 168.000001n V_hig
+ 168.100000n V_hig
+ 168.100001n V_hig
+ 168.200000n V_hig
+ 168.200001n V_hig
+ 168.300000n V_hig
+ 168.300001n V_hig
+ 168.400000n V_hig
+ 168.400001n V_hig
+ 168.500000n V_hig
+ 168.500001n V_hig
+ 168.600000n V_hig
+ 168.600001n V_hig
+ 168.700000n V_hig
+ 168.700001n V_hig
+ 168.800000n V_hig
+ 168.800001n V_hig
+ 168.900000n V_hig
+ 168.900001n V_hig
+ 169.000000n V_hig
+ 169.000001n V_hig
+ 169.100000n V_hig
+ 169.100001n V_hig
+ 169.200000n V_hig
+ 169.200001n V_hig
+ 169.300000n V_hig
+ 169.300001n V_hig
+ 169.400000n V_hig
+ 169.400001n V_hig
+ 169.500000n V_hig
+ 169.500001n V_hig
+ 169.600000n V_hig
+ 169.600001n V_hig
+ 169.700000n V_hig
+ 169.700001n V_hig
+ 169.800000n V_hig
+ 169.800001n V_hig
+ 169.900000n V_hig
+ 169.900001n V_hig
+ 170.000000n V_hig
+ 170.000001n V_low
+ 170.100000n V_low
+ 170.100001n V_low
+ 170.200000n V_low
+ 170.200001n V_low
+ 170.300000n V_low
+ 170.300001n V_low
+ 170.400000n V_low
+ 170.400001n V_low
+ 170.500000n V_low
+ 170.500001n V_low
+ 170.600000n V_low
+ 170.600001n V_low
+ 170.700000n V_low
+ 170.700001n V_low
+ 170.800000n V_low
+ 170.800001n V_low
+ 170.900000n V_low
+ 170.900001n V_low
+ 171.000000n V_low
+ 171.000001n V_hig
+ 171.100000n V_hig
+ 171.100001n V_hig
+ 171.200000n V_hig
+ 171.200001n V_hig
+ 171.300000n V_hig
+ 171.300001n V_hig
+ 171.400000n V_hig
+ 171.400001n V_hig
+ 171.500000n V_hig
+ 171.500001n V_hig
+ 171.600000n V_hig
+ 171.600001n V_hig
+ 171.700000n V_hig
+ 171.700001n V_hig
+ 171.800000n V_hig
+ 171.800001n V_hig
+ 171.900000n V_hig
+ 171.900001n V_hig
+ 172.000000n V_hig
+ 172.000001n V_low
+ 172.100000n V_low
+ 172.100001n V_low
+ 172.200000n V_low
+ 172.200001n V_low
+ 172.300000n V_low
+ 172.300001n V_low
+ 172.400000n V_low
+ 172.400001n V_low
+ 172.500000n V_low
+ 172.500001n V_low
+ 172.600000n V_low
+ 172.600001n V_low
+ 172.700000n V_low
+ 172.700001n V_low
+ 172.800000n V_low
+ 172.800001n V_low
+ 172.900000n V_low
+ 172.900001n V_low
+ 173.000000n V_low
+ 173.000001n V_hig
+ 173.100000n V_hig
+ 173.100001n V_hig
+ 173.200000n V_hig
+ 173.200001n V_hig
+ 173.300000n V_hig
+ 173.300001n V_hig
+ 173.400000n V_hig
+ 173.400001n V_hig
+ 173.500000n V_hig
+ 173.500001n V_hig
+ 173.600000n V_hig
+ 173.600001n V_hig
+ 173.700000n V_hig
+ 173.700001n V_hig
+ 173.800000n V_hig
+ 173.800001n V_hig
+ 173.900000n V_hig
+ 173.900001n V_hig
+ 174.000000n V_hig
+ 174.000001n V_low
+ 174.100000n V_low
+ 174.100001n V_low
+ 174.200000n V_low
+ 174.200001n V_low
+ 174.300000n V_low
+ 174.300001n V_low
+ 174.400000n V_low
+ 174.400001n V_low
+ 174.500000n V_low
+ 174.500001n V_low
+ 174.600000n V_low
+ 174.600001n V_low
+ 174.700000n V_low
+ 174.700001n V_low
+ 174.800000n V_low
+ 174.800001n V_low
+ 174.900000n V_low
+ 174.900001n V_low
+ 175.000000n V_low
+ 175.000001n V_hig
+ 175.100000n V_hig
+ 175.100001n V_hig
+ 175.200000n V_hig
+ 175.200001n V_hig
+ 175.300000n V_hig
+ 175.300001n V_hig
+ 175.400000n V_hig
+ 175.400001n V_hig
+ 175.500000n V_hig
+ 175.500001n V_hig
+ 175.600000n V_hig
+ 175.600001n V_hig
+ 175.700000n V_hig
+ 175.700001n V_hig
+ 175.800000n V_hig
+ 175.800001n V_hig
+ 175.900000n V_hig
+ 175.900001n V_hig
+ 176.000000n V_hig
+ 176.000001n V_hig
+ 176.100000n V_hig
+ 176.100001n V_hig
+ 176.200000n V_hig
+ 176.200001n V_hig
+ 176.300000n V_hig
+ 176.300001n V_hig
+ 176.400000n V_hig
+ 176.400001n V_hig
+ 176.500000n V_hig
+ 176.500001n V_hig
+ 176.600000n V_hig
+ 176.600001n V_hig
+ 176.700000n V_hig
+ 176.700001n V_hig
+ 176.800000n V_hig
+ 176.800001n V_hig
+ 176.900000n V_hig
+ 176.900001n V_hig
+ 177.000000n V_hig
+ 177.000001n V_low
+ 177.100000n V_low
+ 177.100001n V_low
+ 177.200000n V_low
+ 177.200001n V_low
+ 177.300000n V_low
+ 177.300001n V_low
+ 177.400000n V_low
+ 177.400001n V_low
+ 177.500000n V_low
+ 177.500001n V_low
+ 177.600000n V_low
+ 177.600001n V_low
+ 177.700000n V_low
+ 177.700001n V_low
+ 177.800000n V_low
+ 177.800001n V_low
+ 177.900000n V_low
+ 177.900001n V_low
+ 178.000000n V_low
+ 178.000001n V_hig
+ 178.100000n V_hig
+ 178.100001n V_hig
+ 178.200000n V_hig
+ 178.200001n V_hig
+ 178.300000n V_hig
+ 178.300001n V_hig
+ 178.400000n V_hig
+ 178.400001n V_hig
+ 178.500000n V_hig
+ 178.500001n V_hig
+ 178.600000n V_hig
+ 178.600001n V_hig
+ 178.700000n V_hig
+ 178.700001n V_hig
+ 178.800000n V_hig
+ 178.800001n V_hig
+ 178.900000n V_hig
+ 178.900001n V_hig
+ 179.000000n V_hig
+ 179.000001n V_low
+ 179.100000n V_low
+ 179.100001n V_low
+ 179.200000n V_low
+ 179.200001n V_low
+ 179.300000n V_low
+ 179.300001n V_low
+ 179.400000n V_low
+ 179.400001n V_low
+ 179.500000n V_low
+ 179.500001n V_low
+ 179.600000n V_low
+ 179.600001n V_low
+ 179.700000n V_low
+ 179.700001n V_low
+ 179.800000n V_low
+ 179.800001n V_low
+ 179.900000n V_low
+ 179.900001n V_low
+ 180.000000n V_low
+ 180.000001n V_low
+ 180.100000n V_low
+ 180.100001n V_low
+ 180.200000n V_low
+ 180.200001n V_low
+ 180.300000n V_low
+ 180.300001n V_low
+ 180.400000n V_low
+ 180.400001n V_low
+ 180.500000n V_low
+ 180.500001n V_low
+ 180.600000n V_low
+ 180.600001n V_low
+ 180.700000n V_low
+ 180.700001n V_low
+ 180.800000n V_low
+ 180.800001n V_low
+ 180.900000n V_low
+ 180.900001n V_low
+ 181.000000n V_low
+ 181.000001n V_hig
+ 181.100000n V_hig
+ 181.100001n V_hig
+ 181.200000n V_hig
+ 181.200001n V_hig
+ 181.300000n V_hig
+ 181.300001n V_hig
+ 181.400000n V_hig
+ 181.400001n V_hig
+ 181.500000n V_hig
+ 181.500001n V_hig
+ 181.600000n V_hig
+ 181.600001n V_hig
+ 181.700000n V_hig
+ 181.700001n V_hig
+ 181.800000n V_hig
+ 181.800001n V_hig
+ 181.900000n V_hig
+ 181.900001n V_hig
+ 182.000000n V_hig
+ 182.000001n V_low
+ 182.100000n V_low
+ 182.100001n V_low
+ 182.200000n V_low
+ 182.200001n V_low
+ 182.300000n V_low
+ 182.300001n V_low
+ 182.400000n V_low
+ 182.400001n V_low
+ 182.500000n V_low
+ 182.500001n V_low
+ 182.600000n V_low
+ 182.600001n V_low
+ 182.700000n V_low
+ 182.700001n V_low
+ 182.800000n V_low
+ 182.800001n V_low
+ 182.900000n V_low
+ 182.900001n V_low
+ 183.000000n V_low
+ 183.000001n V_low
+ 183.100000n V_low
+ 183.100001n V_low
+ 183.200000n V_low
+ 183.200001n V_low
+ 183.300000n V_low
+ 183.300001n V_low
+ 183.400000n V_low
+ 183.400001n V_low
+ 183.500000n V_low
+ 183.500001n V_low
+ 183.600000n V_low
+ 183.600001n V_low
+ 183.700000n V_low
+ 183.700001n V_low
+ 183.800000n V_low
+ 183.800001n V_low
+ 183.900000n V_low
+ 183.900001n V_low
+ 184.000000n V_low
+ 184.000001n V_low
+ 184.100000n V_low
+ 184.100001n V_low
+ 184.200000n V_low
+ 184.200001n V_low
+ 184.300000n V_low
+ 184.300001n V_low
+ 184.400000n V_low
+ 184.400001n V_low
+ 184.500000n V_low
+ 184.500001n V_low
+ 184.600000n V_low
+ 184.600001n V_low
+ 184.700000n V_low
+ 184.700001n V_low
+ 184.800000n V_low
+ 184.800001n V_low
+ 184.900000n V_low
+ 184.900001n V_low
+ 185.000000n V_low
+ 185.000001n V_low
+ 185.100000n V_low
+ 185.100001n V_low
+ 185.200000n V_low
+ 185.200001n V_low
+ 185.300000n V_low
+ 185.300001n V_low
+ 185.400000n V_low
+ 185.400001n V_low
+ 185.500000n V_low
+ 185.500001n V_low
+ 185.600000n V_low
+ 185.600001n V_low
+ 185.700000n V_low
+ 185.700001n V_low
+ 185.800000n V_low
+ 185.800001n V_low
+ 185.900000n V_low
+ 185.900001n V_low
+ 186.000000n V_low
+ 186.000001n V_hig
+ 186.100000n V_hig
+ 186.100001n V_hig
+ 186.200000n V_hig
+ 186.200001n V_hig
+ 186.300000n V_hig
+ 186.300001n V_hig
+ 186.400000n V_hig
+ 186.400001n V_hig
+ 186.500000n V_hig
+ 186.500001n V_hig
+ 186.600000n V_hig
+ 186.600001n V_hig
+ 186.700000n V_hig
+ 186.700001n V_hig
+ 186.800000n V_hig
+ 186.800001n V_hig
+ 186.900000n V_hig
+ 186.900001n V_hig
+ 187.000000n V_hig
+ 187.000001n V_low
+ 187.100000n V_low
+ 187.100001n V_low
+ 187.200000n V_low
+ 187.200001n V_low
+ 187.300000n V_low
+ 187.300001n V_low
+ 187.400000n V_low
+ 187.400001n V_low
+ 187.500000n V_low
+ 187.500001n V_low
+ 187.600000n V_low
+ 187.600001n V_low
+ 187.700000n V_low
+ 187.700001n V_low
+ 187.800000n V_low
+ 187.800001n V_low
+ 187.900000n V_low
+ 187.900001n V_low
+ 188.000000n V_low
+ 188.000001n V_low
+ 188.100000n V_low
+ 188.100001n V_low
+ 188.200000n V_low
+ 188.200001n V_low
+ 188.300000n V_low
+ 188.300001n V_low
+ 188.400000n V_low
+ 188.400001n V_low
+ 188.500000n V_low
+ 188.500001n V_low
+ 188.600000n V_low
+ 188.600001n V_low
+ 188.700000n V_low
+ 188.700001n V_low
+ 188.800000n V_low
+ 188.800001n V_low
+ 188.900000n V_low
+ 188.900001n V_low
+ 189.000000n V_low
+ 189.000001n V_hig
+ 189.100000n V_hig
+ 189.100001n V_hig
+ 189.200000n V_hig
+ 189.200001n V_hig
+ 189.300000n V_hig
+ 189.300001n V_hig
+ 189.400000n V_hig
+ 189.400001n V_hig
+ 189.500000n V_hig
+ 189.500001n V_hig
+ 189.600000n V_hig
+ 189.600001n V_hig
+ 189.700000n V_hig
+ 189.700001n V_hig
+ 189.800000n V_hig
+ 189.800001n V_hig
+ 189.900000n V_hig
+ 189.900001n V_hig
+ 190.000000n V_hig
+ 190.000001n V_hig
+ 190.100000n V_hig
+ 190.100001n V_hig
+ 190.200000n V_hig
+ 190.200001n V_hig
+ 190.300000n V_hig
+ 190.300001n V_hig
+ 190.400000n V_hig
+ 190.400001n V_hig
+ 190.500000n V_hig
+ 190.500001n V_hig
+ 190.600000n V_hig
+ 190.600001n V_hig
+ 190.700000n V_hig
+ 190.700001n V_hig
+ 190.800000n V_hig
+ 190.800001n V_hig
+ 190.900000n V_hig
+ 190.900001n V_hig
+ 191.000000n V_hig
+ 191.000001n V_hig
+ 191.100000n V_hig
+ 191.100001n V_hig
+ 191.200000n V_hig
+ 191.200001n V_hig
+ 191.300000n V_hig
+ 191.300001n V_hig
+ 191.400000n V_hig
+ 191.400001n V_hig
+ 191.500000n V_hig
+ 191.500001n V_hig
+ 191.600000n V_hig
+ 191.600001n V_hig
+ 191.700000n V_hig
+ 191.700001n V_hig
+ 191.800000n V_hig
+ 191.800001n V_hig
+ 191.900000n V_hig
+ 191.900001n V_hig
+ 192.000000n V_hig
+ 192.000001n V_low
+ 192.100000n V_low
+ 192.100001n V_low
+ 192.200000n V_low
+ 192.200001n V_low
+ 192.300000n V_low
+ 192.300001n V_low
+ 192.400000n V_low
+ 192.400001n V_low
+ 192.500000n V_low
+ 192.500001n V_low
+ 192.600000n V_low
+ 192.600001n V_low
+ 192.700000n V_low
+ 192.700001n V_low
+ 192.800000n V_low
+ 192.800001n V_low
+ 192.900000n V_low
+ 192.900001n V_low
+ 193.000000n V_low
+ 193.000001n V_low
+ 193.100000n V_low
+ 193.100001n V_low
+ 193.200000n V_low
+ 193.200001n V_low
+ 193.300000n V_low
+ 193.300001n V_low
+ 193.400000n V_low
+ 193.400001n V_low
+ 193.500000n V_low
+ 193.500001n V_low
+ 193.600000n V_low
+ 193.600001n V_low
+ 193.700000n V_low
+ 193.700001n V_low
+ 193.800000n V_low
+ 193.800001n V_low
+ 193.900000n V_low
+ 193.900001n V_low
+ 194.000000n V_low
+ 194.000001n V_low
+ 194.100000n V_low
+ 194.100001n V_low
+ 194.200000n V_low
+ 194.200001n V_low
+ 194.300000n V_low
+ 194.300001n V_low
+ 194.400000n V_low
+ 194.400001n V_low
+ 194.500000n V_low
+ 194.500001n V_low
+ 194.600000n V_low
+ 194.600001n V_low
+ 194.700000n V_low
+ 194.700001n V_low
+ 194.800000n V_low
+ 194.800001n V_low
+ 194.900000n V_low
+ 194.900001n V_low
+ 195.000000n V_low
+ 195.000001n V_low
+ 195.100000n V_low
+ 195.100001n V_low
+ 195.200000n V_low
+ 195.200001n V_low
+ 195.300000n V_low
+ 195.300001n V_low
+ 195.400000n V_low
+ 195.400001n V_low
+ 195.500000n V_low
+ 195.500001n V_low
+ 195.600000n V_low
+ 195.600001n V_low
+ 195.700000n V_low
+ 195.700001n V_low
+ 195.800000n V_low
+ 195.800001n V_low
+ 195.900000n V_low
+ 195.900001n V_low
+ 196.000000n V_low
+ 196.000001n V_hig
+ 196.100000n V_hig
+ 196.100001n V_hig
+ 196.200000n V_hig
+ 196.200001n V_hig
+ 196.300000n V_hig
+ 196.300001n V_hig
+ 196.400000n V_hig
+ 196.400001n V_hig
+ 196.500000n V_hig
+ 196.500001n V_hig
+ 196.600000n V_hig
+ 196.600001n V_hig
+ 196.700000n V_hig
+ 196.700001n V_hig
+ 196.800000n V_hig
+ 196.800001n V_hig
+ 196.900000n V_hig
+ 196.900001n V_hig
+ 197.000000n V_hig
+ 197.000001n V_hig
+ 197.100000n V_hig
+ 197.100001n V_hig
+ 197.200000n V_hig
+ 197.200001n V_hig
+ 197.300000n V_hig
+ 197.300001n V_hig
+ 197.400000n V_hig
+ 197.400001n V_hig
+ 197.500000n V_hig
+ 197.500001n V_hig
+ 197.600000n V_hig
+ 197.600001n V_hig
+ 197.700000n V_hig
+ 197.700001n V_hig
+ 197.800000n V_hig
+ 197.800001n V_hig
+ 197.900000n V_hig
+ 197.900001n V_hig
+ 198.000000n V_hig
+ 198.000001n V_hig
+ 198.100000n V_hig
+ 198.100001n V_hig
+ 198.200000n V_hig
+ 198.200001n V_hig
+ 198.300000n V_hig
+ 198.300001n V_hig
+ 198.400000n V_hig
+ 198.400001n V_hig
+ 198.500000n V_hig
+ 198.500001n V_hig
+ 198.600000n V_hig
+ 198.600001n V_hig
+ 198.700000n V_hig
+ 198.700001n V_hig
+ 198.800000n V_hig
+ 198.800001n V_hig
+ 198.900000n V_hig
+ 198.900001n V_hig
+ 199.000000n V_hig
+ 199.000001n V_low
+ 199.100000n V_low
+ 199.100001n V_low
+ 199.200000n V_low
+ 199.200001n V_low
+ 199.300000n V_low
+ 199.300001n V_low
+ 199.400000n V_low
+ 199.400001n V_low
+ 199.500000n V_low
+ 199.500001n V_low
+ 199.600000n V_low
+ 199.600001n V_low
+ 199.700000n V_low
+ 199.700001n V_low
+ 199.800000n V_low
+ 199.800001n V_low
+ 199.900000n V_low
+ 199.900001n V_low
+ 200.000000n V_low
+ 200.000001n V_low
+ 200.100000n V_low
+ 200.100001n V_low
+ 200.200000n V_low
+ 200.200001n V_low
+ 200.300000n V_low
+ 200.300001n V_low
+ 200.400000n V_low
+ 200.400001n V_low
+ 200.500000n V_low
+ 200.500001n V_low
+ 200.600000n V_low
+ 200.600001n V_low
+ 200.700000n V_low
+ 200.700001n V_low
+ 200.800000n V_low
+ 200.800001n V_low
+ 200.900000n V_low
+ 200.900001n V_low
+ 201.000000n V_low
+ 201.000001n V_low
+ 201.100000n V_low
+ 201.100001n V_low
+ 201.200000n V_low
+ 201.200001n V_low
+ 201.300000n V_low
+ 201.300001n V_low
+ 201.400000n V_low
+ 201.400001n V_low
+ 201.500000n V_low
+ 201.500001n V_low
+ 201.600000n V_low
+ 201.600001n V_low
+ 201.700000n V_low
+ 201.700001n V_low
+ 201.800000n V_low
+ 201.800001n V_low
+ 201.900000n V_low
+ 201.900001n V_low
+ 202.000000n V_low
+ 202.000001n V_low
+ 202.100000n V_low
+ 202.100001n V_low
+ 202.200000n V_low
+ 202.200001n V_low
+ 202.300000n V_low
+ 202.300001n V_low
+ 202.400000n V_low
+ 202.400001n V_low
+ 202.500000n V_low
+ 202.500001n V_low
+ 202.600000n V_low
+ 202.600001n V_low
+ 202.700000n V_low
+ 202.700001n V_low
+ 202.800000n V_low
+ 202.800001n V_low
+ 202.900000n V_low
+ 202.900001n V_low
+ 203.000000n V_low
+ 203.000001n V_low
+ 203.100000n V_low
+ 203.100001n V_low
+ 203.200000n V_low
+ 203.200001n V_low
+ 203.300000n V_low
+ 203.300001n V_low
+ 203.400000n V_low
+ 203.400001n V_low
+ 203.500000n V_low
+ 203.500001n V_low
+ 203.600000n V_low
+ 203.600001n V_low
+ 203.700000n V_low
+ 203.700001n V_low
+ 203.800000n V_low
+ 203.800001n V_low
+ 203.900000n V_low
+ 203.900001n V_low
+ 204.000000n V_low
+ 204.000001n V_hig
+ 204.100000n V_hig
+ 204.100001n V_hig
+ 204.200000n V_hig
+ 204.200001n V_hig
+ 204.300000n V_hig
+ 204.300001n V_hig
+ 204.400000n V_hig
+ 204.400001n V_hig
+ 204.500000n V_hig
+ 204.500001n V_hig
+ 204.600000n V_hig
+ 204.600001n V_hig
+ 204.700000n V_hig
+ 204.700001n V_hig
+ 204.800000n V_hig
+ 204.800001n V_hig
+ 204.900000n V_hig
+ 204.900001n V_hig
+ 205.000000n V_hig
+ 205.000001n V_low
+ 205.100000n V_low
+ 205.100001n V_low
+ 205.200000n V_low
+ 205.200001n V_low
+ 205.300000n V_low
+ 205.300001n V_low
+ 205.400000n V_low
+ 205.400001n V_low
+ 205.500000n V_low
+ 205.500001n V_low
+ 205.600000n V_low
+ 205.600001n V_low
+ 205.700000n V_low
+ 205.700001n V_low
+ 205.800000n V_low
+ 205.800001n V_low
+ 205.900000n V_low
+ 205.900001n V_low
+ 206.000000n V_low
+ 206.000001n V_low
+ 206.100000n V_low
+ 206.100001n V_low
+ 206.200000n V_low
+ 206.200001n V_low
+ 206.300000n V_low
+ 206.300001n V_low
+ 206.400000n V_low
+ 206.400001n V_low
+ 206.500000n V_low
+ 206.500001n V_low
+ 206.600000n V_low
+ 206.600001n V_low
+ 206.700000n V_low
+ 206.700001n V_low
+ 206.800000n V_low
+ 206.800001n V_low
+ 206.900000n V_low
+ 206.900001n V_low
+ 207.000000n V_low
+ 207.000001n V_low
+ 207.100000n V_low
+ 207.100001n V_low
+ 207.200000n V_low
+ 207.200001n V_low
+ 207.300000n V_low
+ 207.300001n V_low
+ 207.400000n V_low
+ 207.400001n V_low
+ 207.500000n V_low
+ 207.500001n V_low
+ 207.600000n V_low
+ 207.600001n V_low
+ 207.700000n V_low
+ 207.700001n V_low
+ 207.800000n V_low
+ 207.800001n V_low
+ 207.900000n V_low
+ 207.900001n V_low
+ 208.000000n V_low
+ 208.000001n V_low
+ 208.100000n V_low
+ 208.100001n V_low
+ 208.200000n V_low
+ 208.200001n V_low
+ 208.300000n V_low
+ 208.300001n V_low
+ 208.400000n V_low
+ 208.400001n V_low
+ 208.500000n V_low
+ 208.500001n V_low
+ 208.600000n V_low
+ 208.600001n V_low
+ 208.700000n V_low
+ 208.700001n V_low
+ 208.800000n V_low
+ 208.800001n V_low
+ 208.900000n V_low
+ 208.900001n V_low
+ 209.000000n V_low
+ 209.000001n V_hig
+ 209.100000n V_hig
+ 209.100001n V_hig
+ 209.200000n V_hig
+ 209.200001n V_hig
+ 209.300000n V_hig
+ 209.300001n V_hig
+ 209.400000n V_hig
+ 209.400001n V_hig
+ 209.500000n V_hig
+ 209.500001n V_hig
+ 209.600000n V_hig
+ 209.600001n V_hig
+ 209.700000n V_hig
+ 209.700001n V_hig
+ 209.800000n V_hig
+ 209.800001n V_hig
+ 209.900000n V_hig
+ 209.900001n V_hig
+ 210.000000n V_hig
+ 210.000001n V_hig
+ 210.100000n V_hig
+ 210.100001n V_hig
+ 210.200000n V_hig
+ 210.200001n V_hig
+ 210.300000n V_hig
+ 210.300001n V_hig
+ 210.400000n V_hig
+ 210.400001n V_hig
+ 210.500000n V_hig
+ 210.500001n V_hig
+ 210.600000n V_hig
+ 210.600001n V_hig
+ 210.700000n V_hig
+ 210.700001n V_hig
+ 210.800000n V_hig
+ 210.800001n V_hig
+ 210.900000n V_hig
+ 210.900001n V_hig
+ 211.000000n V_hig
+ 211.000001n V_low
+ 211.100000n V_low
+ 211.100001n V_low
+ 211.200000n V_low
+ 211.200001n V_low
+ 211.300000n V_low
+ 211.300001n V_low
+ 211.400000n V_low
+ 211.400001n V_low
+ 211.500000n V_low
+ 211.500001n V_low
+ 211.600000n V_low
+ 211.600001n V_low
+ 211.700000n V_low
+ 211.700001n V_low
+ 211.800000n V_low
+ 211.800001n V_low
+ 211.900000n V_low
+ 211.900001n V_low
+ 212.000000n V_low
+ 212.000001n V_hig
+ 212.100000n V_hig
+ 212.100001n V_hig
+ 212.200000n V_hig
+ 212.200001n V_hig
+ 212.300000n V_hig
+ 212.300001n V_hig
+ 212.400000n V_hig
+ 212.400001n V_hig
+ 212.500000n V_hig
+ 212.500001n V_hig
+ 212.600000n V_hig
+ 212.600001n V_hig
+ 212.700000n V_hig
+ 212.700001n V_hig
+ 212.800000n V_hig
+ 212.800001n V_hig
+ 212.900000n V_hig
+ 212.900001n V_hig
+ 213.000000n V_hig
+ 213.000001n V_hig
+ 213.100000n V_hig
+ 213.100001n V_hig
+ 213.200000n V_hig
+ 213.200001n V_hig
+ 213.300000n V_hig
+ 213.300001n V_hig
+ 213.400000n V_hig
+ 213.400001n V_hig
+ 213.500000n V_hig
+ 213.500001n V_hig
+ 213.600000n V_hig
+ 213.600001n V_hig
+ 213.700000n V_hig
+ 213.700001n V_hig
+ 213.800000n V_hig
+ 213.800001n V_hig
+ 213.900000n V_hig
+ 213.900001n V_hig
+ 214.000000n V_hig
+ 214.000001n V_hig
+ 214.100000n V_hig
+ 214.100001n V_hig
+ 214.200000n V_hig
+ 214.200001n V_hig
+ 214.300000n V_hig
+ 214.300001n V_hig
+ 214.400000n V_hig
+ 214.400001n V_hig
+ 214.500000n V_hig
+ 214.500001n V_hig
+ 214.600000n V_hig
+ 214.600001n V_hig
+ 214.700000n V_hig
+ 214.700001n V_hig
+ 214.800000n V_hig
+ 214.800001n V_hig
+ 214.900000n V_hig
+ 214.900001n V_hig
+ 215.000000n V_hig
+ 215.000001n V_hig
+ 215.100000n V_hig
+ 215.100001n V_hig
+ 215.200000n V_hig
+ 215.200001n V_hig
+ 215.300000n V_hig
+ 215.300001n V_hig
+ 215.400000n V_hig
+ 215.400001n V_hig
+ 215.500000n V_hig
+ 215.500001n V_hig
+ 215.600000n V_hig
+ 215.600001n V_hig
+ 215.700000n V_hig
+ 215.700001n V_hig
+ 215.800000n V_hig
+ 215.800001n V_hig
+ 215.900000n V_hig
+ 215.900001n V_hig
+ 216.000000n V_hig
+ 216.000001n V_low
+ 216.100000n V_low
+ 216.100001n V_low
+ 216.200000n V_low
+ 216.200001n V_low
+ 216.300000n V_low
+ 216.300001n V_low
+ 216.400000n V_low
+ 216.400001n V_low
+ 216.500000n V_low
+ 216.500001n V_low
+ 216.600000n V_low
+ 216.600001n V_low
+ 216.700000n V_low
+ 216.700001n V_low
+ 216.800000n V_low
+ 216.800001n V_low
+ 216.900000n V_low
+ 216.900001n V_low
+ 217.000000n V_low
+ 217.000001n V_low
+ 217.100000n V_low
+ 217.100001n V_low
+ 217.200000n V_low
+ 217.200001n V_low
+ 217.300000n V_low
+ 217.300001n V_low
+ 217.400000n V_low
+ 217.400001n V_low
+ 217.500000n V_low
+ 217.500001n V_low
+ 217.600000n V_low
+ 217.600001n V_low
+ 217.700000n V_low
+ 217.700001n V_low
+ 217.800000n V_low
+ 217.800001n V_low
+ 217.900000n V_low
+ 217.900001n V_low
+ 218.000000n V_low
+ 218.000001n V_hig
+ 218.100000n V_hig
+ 218.100001n V_hig
+ 218.200000n V_hig
+ 218.200001n V_hig
+ 218.300000n V_hig
+ 218.300001n V_hig
+ 218.400000n V_hig
+ 218.400001n V_hig
+ 218.500000n V_hig
+ 218.500001n V_hig
+ 218.600000n V_hig
+ 218.600001n V_hig
+ 218.700000n V_hig
+ 218.700001n V_hig
+ 218.800000n V_hig
+ 218.800001n V_hig
+ 218.900000n V_hig
+ 218.900001n V_hig
+ 219.000000n V_hig
+ 219.000001n V_low
+ 219.100000n V_low
+ 219.100001n V_low
+ 219.200000n V_low
+ 219.200001n V_low
+ 219.300000n V_low
+ 219.300001n V_low
+ 219.400000n V_low
+ 219.400001n V_low
+ 219.500000n V_low
+ 219.500001n V_low
+ 219.600000n V_low
+ 219.600001n V_low
+ 219.700000n V_low
+ 219.700001n V_low
+ 219.800000n V_low
+ 219.800001n V_low
+ 219.900000n V_low
+ 219.900001n V_low
+ 220.000000n V_low
+ 220.000001n V_low
+ 220.100000n V_low
+ 220.100001n V_low
+ 220.200000n V_low
+ 220.200001n V_low
+ 220.300000n V_low
+ 220.300001n V_low
+ 220.400000n V_low
+ 220.400001n V_low
+ 220.500000n V_low
+ 220.500001n V_low
+ 220.600000n V_low
+ 220.600001n V_low
+ 220.700000n V_low
+ 220.700001n V_low
+ 220.800000n V_low
+ 220.800001n V_low
+ 220.900000n V_low
+ 220.900001n V_low
+ 221.000000n V_low
+ 221.000001n V_hig
+ 221.100000n V_hig
+ 221.100001n V_hig
+ 221.200000n V_hig
+ 221.200001n V_hig
+ 221.300000n V_hig
+ 221.300001n V_hig
+ 221.400000n V_hig
+ 221.400001n V_hig
+ 221.500000n V_hig
+ 221.500001n V_hig
+ 221.600000n V_hig
+ 221.600001n V_hig
+ 221.700000n V_hig
+ 221.700001n V_hig
+ 221.800000n V_hig
+ 221.800001n V_hig
+ 221.900000n V_hig
+ 221.900001n V_hig
+ 222.000000n V_hig
+ 222.000001n V_hig
+ 222.100000n V_hig
+ 222.100001n V_hig
+ 222.200000n V_hig
+ 222.200001n V_hig
+ 222.300000n V_hig
+ 222.300001n V_hig
+ 222.400000n V_hig
+ 222.400001n V_hig
+ 222.500000n V_hig
+ 222.500001n V_hig
+ 222.600000n V_hig
+ 222.600001n V_hig
+ 222.700000n V_hig
+ 222.700001n V_hig
+ 222.800000n V_hig
+ 222.800001n V_hig
+ 222.900000n V_hig
+ 222.900001n V_hig
+ 223.000000n V_hig
+ 223.000001n V_low
+ 223.100000n V_low
+ 223.100001n V_low
+ 223.200000n V_low
+ 223.200001n V_low
+ 223.300000n V_low
+ 223.300001n V_low
+ 223.400000n V_low
+ 223.400001n V_low
+ 223.500000n V_low
+ 223.500001n V_low
+ 223.600000n V_low
+ 223.600001n V_low
+ 223.700000n V_low
+ 223.700001n V_low
+ 223.800000n V_low
+ 223.800001n V_low
+ 223.900000n V_low
+ 223.900001n V_low
+ 224.000000n V_low
+ 224.000001n V_low
+ 224.100000n V_low
+ 224.100001n V_low
+ 224.200000n V_low
+ 224.200001n V_low
+ 224.300000n V_low
+ 224.300001n V_low
+ 224.400000n V_low
+ 224.400001n V_low
+ 224.500000n V_low
+ 224.500001n V_low
+ 224.600000n V_low
+ 224.600001n V_low
+ 224.700000n V_low
+ 224.700001n V_low
+ 224.800000n V_low
+ 224.800001n V_low
+ 224.900000n V_low
+ 224.900001n V_low
+ 225.000000n V_low
+ 225.000001n V_low
+ 225.100000n V_low
+ 225.100001n V_low
+ 225.200000n V_low
+ 225.200001n V_low
+ 225.300000n V_low
+ 225.300001n V_low
+ 225.400000n V_low
+ 225.400001n V_low
+ 225.500000n V_low
+ 225.500001n V_low
+ 225.600000n V_low
+ 225.600001n V_low
+ 225.700000n V_low
+ 225.700001n V_low
+ 225.800000n V_low
+ 225.800001n V_low
+ 225.900000n V_low
+ 225.900001n V_low
+ 226.000000n V_low
+ 226.000001n V_low
+ 226.100000n V_low
+ 226.100001n V_low
+ 226.200000n V_low
+ 226.200001n V_low
+ 226.300000n V_low
+ 226.300001n V_low
+ 226.400000n V_low
+ 226.400001n V_low
+ 226.500000n V_low
+ 226.500001n V_low
+ 226.600000n V_low
+ 226.600001n V_low
+ 226.700000n V_low
+ 226.700001n V_low
+ 226.800000n V_low
+ 226.800001n V_low
+ 226.900000n V_low
+ 226.900001n V_low
+ 227.000000n V_low
+ 227.000001n V_hig
+ 227.100000n V_hig
+ 227.100001n V_hig
+ 227.200000n V_hig
+ 227.200001n V_hig
+ 227.300000n V_hig
+ 227.300001n V_hig
+ 227.400000n V_hig
+ 227.400001n V_hig
+ 227.500000n V_hig
+ 227.500001n V_hig
+ 227.600000n V_hig
+ 227.600001n V_hig
+ 227.700000n V_hig
+ 227.700001n V_hig
+ 227.800000n V_hig
+ 227.800001n V_hig
+ 227.900000n V_hig
+ 227.900001n V_hig
+ 228.000000n V_hig
+ 228.000001n V_low
+ 228.100000n V_low
+ 228.100001n V_low
+ 228.200000n V_low
+ 228.200001n V_low
+ 228.300000n V_low
+ 228.300001n V_low
+ 228.400000n V_low
+ 228.400001n V_low
+ 228.500000n V_low
+ 228.500001n V_low
+ 228.600000n V_low
+ 228.600001n V_low
+ 228.700000n V_low
+ 228.700001n V_low
+ 228.800000n V_low
+ 228.800001n V_low
+ 228.900000n V_low
+ 228.900001n V_low
+ 229.000000n V_low
+ 229.000001n V_hig
+ 229.100000n V_hig
+ 229.100001n V_hig
+ 229.200000n V_hig
+ 229.200001n V_hig
+ 229.300000n V_hig
+ 229.300001n V_hig
+ 229.400000n V_hig
+ 229.400001n V_hig
+ 229.500000n V_hig
+ 229.500001n V_hig
+ 229.600000n V_hig
+ 229.600001n V_hig
+ 229.700000n V_hig
+ 229.700001n V_hig
+ 229.800000n V_hig
+ 229.800001n V_hig
+ 229.900000n V_hig
+ 229.900001n V_hig
+ 230.000000n V_hig
+ 230.000001n V_hig
+ 230.100000n V_hig
+ 230.100001n V_hig
+ 230.200000n V_hig
+ 230.200001n V_hig
+ 230.300000n V_hig
+ 230.300001n V_hig
+ 230.400000n V_hig
+ 230.400001n V_hig
+ 230.500000n V_hig
+ 230.500001n V_hig
+ 230.600000n V_hig
+ 230.600001n V_hig
+ 230.700000n V_hig
+ 230.700001n V_hig
+ 230.800000n V_hig
+ 230.800001n V_hig
+ 230.900000n V_hig
+ 230.900001n V_hig
+ 231.000000n V_hig
+ 231.000001n V_hig
+ 231.100000n V_hig
+ 231.100001n V_hig
+ 231.200000n V_hig
+ 231.200001n V_hig
+ 231.300000n V_hig
+ 231.300001n V_hig
+ 231.400000n V_hig
+ 231.400001n V_hig
+ 231.500000n V_hig
+ 231.500001n V_hig
+ 231.600000n V_hig
+ 231.600001n V_hig
+ 231.700000n V_hig
+ 231.700001n V_hig
+ 231.800000n V_hig
+ 231.800001n V_hig
+ 231.900000n V_hig
+ 231.900001n V_hig
+ 232.000000n V_hig
+ 232.000001n V_hig
+ 232.100000n V_hig
+ 232.100001n V_hig
+ 232.200000n V_hig
+ 232.200001n V_hig
+ 232.300000n V_hig
+ 232.300001n V_hig
+ 232.400000n V_hig
+ 232.400001n V_hig
+ 232.500000n V_hig
+ 232.500001n V_hig
+ 232.600000n V_hig
+ 232.600001n V_hig
+ 232.700000n V_hig
+ 232.700001n V_hig
+ 232.800000n V_hig
+ 232.800001n V_hig
+ 232.900000n V_hig
+ 232.900001n V_hig
+ 233.000000n V_hig
+ 233.000001n V_hig
+ 233.100000n V_hig
+ 233.100001n V_hig
+ 233.200000n V_hig
+ 233.200001n V_hig
+ 233.300000n V_hig
+ 233.300001n V_hig
+ 233.400000n V_hig
+ 233.400001n V_hig
+ 233.500000n V_hig
+ 233.500001n V_hig
+ 233.600000n V_hig
+ 233.600001n V_hig
+ 233.700000n V_hig
+ 233.700001n V_hig
+ 233.800000n V_hig
+ 233.800001n V_hig
+ 233.900000n V_hig
+ 233.900001n V_hig
+ 234.000000n V_hig
+ 234.000001n V_hig
+ 234.100000n V_hig
+ 234.100001n V_hig
+ 234.200000n V_hig
+ 234.200001n V_hig
+ 234.300000n V_hig
+ 234.300001n V_hig
+ 234.400000n V_hig
+ 234.400001n V_hig
+ 234.500000n V_hig
+ 234.500001n V_hig
+ 234.600000n V_hig
+ 234.600001n V_hig
+ 234.700000n V_hig
+ 234.700001n V_hig
+ 234.800000n V_hig
+ 234.800001n V_hig
+ 234.900000n V_hig
+ 234.900001n V_hig
+ 235.000000n V_hig
+ 235.000001n V_hig
+ 235.100000n V_hig
+ 235.100001n V_hig
+ 235.200000n V_hig
+ 235.200001n V_hig
+ 235.300000n V_hig
+ 235.300001n V_hig
+ 235.400000n V_hig
+ 235.400001n V_hig
+ 235.500000n V_hig
+ 235.500001n V_hig
+ 235.600000n V_hig
+ 235.600001n V_hig
+ 235.700000n V_hig
+ 235.700001n V_hig
+ 235.800000n V_hig
+ 235.800001n V_hig
+ 235.900000n V_hig
+ 235.900001n V_hig
+ 236.000000n V_hig
+ 236.000001n V_hig
+ 236.100000n V_hig
+ 236.100001n V_hig
+ 236.200000n V_hig
+ 236.200001n V_hig
+ 236.300000n V_hig
+ 236.300001n V_hig
+ 236.400000n V_hig
+ 236.400001n V_hig
+ 236.500000n V_hig
+ 236.500001n V_hig
+ 236.600000n V_hig
+ 236.600001n V_hig
+ 236.700000n V_hig
+ 236.700001n V_hig
+ 236.800000n V_hig
+ 236.800001n V_hig
+ 236.900000n V_hig
+ 236.900001n V_hig
+ 237.000000n V_hig
+ 237.000001n V_low
+ 237.100000n V_low
+ 237.100001n V_low
+ 237.200000n V_low
+ 237.200001n V_low
+ 237.300000n V_low
+ 237.300001n V_low
+ 237.400000n V_low
+ 237.400001n V_low
+ 237.500000n V_low
+ 237.500001n V_low
+ 237.600000n V_low
+ 237.600001n V_low
+ 237.700000n V_low
+ 237.700001n V_low
+ 237.800000n V_low
+ 237.800001n V_low
+ 237.900000n V_low
+ 237.900001n V_low
+ 238.000000n V_low
+ 238.000001n V_hig
+ 238.100000n V_hig
+ 238.100001n V_hig
+ 238.200000n V_hig
+ 238.200001n V_hig
+ 238.300000n V_hig
+ 238.300001n V_hig
+ 238.400000n V_hig
+ 238.400001n V_hig
+ 238.500000n V_hig
+ 238.500001n V_hig
+ 238.600000n V_hig
+ 238.600001n V_hig
+ 238.700000n V_hig
+ 238.700001n V_hig
+ 238.800000n V_hig
+ 238.800001n V_hig
+ 238.900000n V_hig
+ 238.900001n V_hig
+ 239.000000n V_hig
+ 239.000001n V_low
+ 239.100000n V_low
+ 239.100001n V_low
+ 239.200000n V_low
+ 239.200001n V_low
+ 239.300000n V_low
+ 239.300001n V_low
+ 239.400000n V_low
+ 239.400001n V_low
+ 239.500000n V_low
+ 239.500001n V_low
+ 239.600000n V_low
+ 239.600001n V_low
+ 239.700000n V_low
+ 239.700001n V_low
+ 239.800000n V_low
+ 239.800001n V_low
+ 239.900000n V_low
+ 239.900001n V_low
+ 240.000000n V_low
+ 240.000001n V_low
+ 240.100000n V_low
+ 240.100001n V_low
+ 240.200000n V_low
+ 240.200001n V_low
+ 240.300000n V_low
+ 240.300001n V_low
+ 240.400000n V_low
+ 240.400001n V_low
+ 240.500000n V_low
+ 240.500001n V_low
+ 240.600000n V_low
+ 240.600001n V_low
+ 240.700000n V_low
+ 240.700001n V_low
+ 240.800000n V_low
+ 240.800001n V_low
+ 240.900000n V_low
+ 240.900001n V_low
+ 241.000000n V_low
+ 241.000001n V_hig
+ 241.100000n V_hig
+ 241.100001n V_hig
+ 241.200000n V_hig
+ 241.200001n V_hig
+ 241.300000n V_hig
+ 241.300001n V_hig
+ 241.400000n V_hig
+ 241.400001n V_hig
+ 241.500000n V_hig
+ 241.500001n V_hig
+ 241.600000n V_hig
+ 241.600001n V_hig
+ 241.700000n V_hig
+ 241.700001n V_hig
+ 241.800000n V_hig
+ 241.800001n V_hig
+ 241.900000n V_hig
+ 241.900001n V_hig
+ 242.000000n V_hig
+ 242.000001n V_low
+ 242.100000n V_low
+ 242.100001n V_low
+ 242.200000n V_low
+ 242.200001n V_low
+ 242.300000n V_low
+ 242.300001n V_low
+ 242.400000n V_low
+ 242.400001n V_low
+ 242.500000n V_low
+ 242.500001n V_low
+ 242.600000n V_low
+ 242.600001n V_low
+ 242.700000n V_low
+ 242.700001n V_low
+ 242.800000n V_low
+ 242.800001n V_low
+ 242.900000n V_low
+ 242.900001n V_low
+ 243.000000n V_low
+ 243.000001n V_hig
+ 243.100000n V_hig
+ 243.100001n V_hig
+ 243.200000n V_hig
+ 243.200001n V_hig
+ 243.300000n V_hig
+ 243.300001n V_hig
+ 243.400000n V_hig
+ 243.400001n V_hig
+ 243.500000n V_hig
+ 243.500001n V_hig
+ 243.600000n V_hig
+ 243.600001n V_hig
+ 243.700000n V_hig
+ 243.700001n V_hig
+ 243.800000n V_hig
+ 243.800001n V_hig
+ 243.900000n V_hig
+ 243.900001n V_hig
+ 244.000000n V_hig
+ 244.000001n V_hig
+ 244.100000n V_hig
+ 244.100001n V_hig
+ 244.200000n V_hig
+ 244.200001n V_hig
+ 244.300000n V_hig
+ 244.300001n V_hig
+ 244.400000n V_hig
+ 244.400001n V_hig
+ 244.500000n V_hig
+ 244.500001n V_hig
+ 244.600000n V_hig
+ 244.600001n V_hig
+ 244.700000n V_hig
+ 244.700001n V_hig
+ 244.800000n V_hig
+ 244.800001n V_hig
+ 244.900000n V_hig
+ 244.900001n V_hig
+ 245.000000n V_hig
+ 245.000001n V_low
+ 245.100000n V_low
+ 245.100001n V_low
+ 245.200000n V_low
+ 245.200001n V_low
+ 245.300000n V_low
+ 245.300001n V_low
+ 245.400000n V_low
+ 245.400001n V_low
+ 245.500000n V_low
+ 245.500001n V_low
+ 245.600000n V_low
+ 245.600001n V_low
+ 245.700000n V_low
+ 245.700001n V_low
+ 245.800000n V_low
+ 245.800001n V_low
+ 245.900000n V_low
+ 245.900001n V_low
+ 246.000000n V_low
+ 246.000001n V_hig
+ 246.100000n V_hig
+ 246.100001n V_hig
+ 246.200000n V_hig
+ 246.200001n V_hig
+ 246.300000n V_hig
+ 246.300001n V_hig
+ 246.400000n V_hig
+ 246.400001n V_hig
+ 246.500000n V_hig
+ 246.500001n V_hig
+ 246.600000n V_hig
+ 246.600001n V_hig
+ 246.700000n V_hig
+ 246.700001n V_hig
+ 246.800000n V_hig
+ 246.800001n V_hig
+ 246.900000n V_hig
+ 246.900001n V_hig
+ 247.000000n V_hig
+ 247.000001n V_hig
+ 247.100000n V_hig
+ 247.100001n V_hig
+ 247.200000n V_hig
+ 247.200001n V_hig
+ 247.300000n V_hig
+ 247.300001n V_hig
+ 247.400000n V_hig
+ 247.400001n V_hig
+ 247.500000n V_hig
+ 247.500001n V_hig
+ 247.600000n V_hig
+ 247.600001n V_hig
+ 247.700000n V_hig
+ 247.700001n V_hig
+ 247.800000n V_hig
+ 247.800001n V_hig
+ 247.900000n V_hig
+ 247.900001n V_hig
+ 248.000000n V_hig
+ 248.000001n V_hig
+ 248.100000n V_hig
+ 248.100001n V_hig
+ 248.200000n V_hig
+ 248.200001n V_hig
+ 248.300000n V_hig
+ 248.300001n V_hig
+ 248.400000n V_hig
+ 248.400001n V_hig
+ 248.500000n V_hig
+ 248.500001n V_hig
+ 248.600000n V_hig
+ 248.600001n V_hig
+ 248.700000n V_hig
+ 248.700001n V_hig
+ 248.800000n V_hig
+ 248.800001n V_hig
+ 248.900000n V_hig
+ 248.900001n V_hig
+ 249.000000n V_hig
+ 249.000001n V_low
+ 249.100000n V_low
+ 249.100001n V_low
+ 249.200000n V_low
+ 249.200001n V_low
+ 249.300000n V_low
+ 249.300001n V_low
+ 249.400000n V_low
+ 249.400001n V_low
+ 249.500000n V_low
+ 249.500001n V_low
+ 249.600000n V_low
+ 249.600001n V_low
+ 249.700000n V_low
+ 249.700001n V_low
+ 249.800000n V_low
+ 249.800001n V_low
+ 249.900000n V_low
+ 249.900001n V_low
+ 250.000000n V_low
+ 250.000001n V_low
+ 250.100000n V_low
+ 250.100001n V_low
+ 250.200000n V_low
+ 250.200001n V_low
+ 250.300000n V_low
+ 250.300001n V_low
+ 250.400000n V_low
+ 250.400001n V_low
+ 250.500000n V_low
+ 250.500001n V_low
+ 250.600000n V_low
+ 250.600001n V_low
+ 250.700000n V_low
+ 250.700001n V_low
+ 250.800000n V_low
+ 250.800001n V_low
+ 250.900000n V_low
+ 250.900001n V_low
+ 251.000000n V_low
+ 251.000001n V_low
+ 251.100000n V_low
+ 251.100001n V_low
+ 251.200000n V_low
+ 251.200001n V_low
+ 251.300000n V_low
+ 251.300001n V_low
+ 251.400000n V_low
+ 251.400001n V_low
+ 251.500000n V_low
+ 251.500001n V_low
+ 251.600000n V_low
+ 251.600001n V_low
+ 251.700000n V_low
+ 251.700001n V_low
+ 251.800000n V_low
+ 251.800001n V_low
+ 251.900000n V_low
+ 251.900001n V_low
+ 252.000000n V_low
+ 252.000001n V_low
+ 252.100000n V_low
+ 252.100001n V_low
+ 252.200000n V_low
+ 252.200001n V_low
+ 252.300000n V_low
+ 252.300001n V_low
+ 252.400000n V_low
+ 252.400001n V_low
+ 252.500000n V_low
+ 252.500001n V_low
+ 252.600000n V_low
+ 252.600001n V_low
+ 252.700000n V_low
+ 252.700001n V_low
+ 252.800000n V_low
+ 252.800001n V_low
+ 252.900000n V_low
+ 252.900001n V_low
+ 253.000000n V_low
+ 253.000001n V_hig
+ 253.100000n V_hig
+ 253.100001n V_hig
+ 253.200000n V_hig
+ 253.200001n V_hig
+ 253.300000n V_hig
+ 253.300001n V_hig
+ 253.400000n V_hig
+ 253.400001n V_hig
+ 253.500000n V_hig
+ 253.500001n V_hig
+ 253.600000n V_hig
+ 253.600001n V_hig
+ 253.700000n V_hig
+ 253.700001n V_hig
+ 253.800000n V_hig
+ 253.800001n V_hig
+ 253.900000n V_hig
+ 253.900001n V_hig
+ 254.000000n V_hig
+ 254.000001n V_low
+ 254.100000n V_low
+ 254.100001n V_low
+ 254.200000n V_low
+ 254.200001n V_low
+ 254.300000n V_low
+ 254.300001n V_low
+ 254.400000n V_low
+ 254.400001n V_low
+ 254.500000n V_low
+ 254.500001n V_low
+ 254.600000n V_low
+ 254.600001n V_low
+ 254.700000n V_low
+ 254.700001n V_low
+ 254.800000n V_low
+ 254.800001n V_low
+ 254.900000n V_low
+ 254.900001n V_low
+ 255.000000n V_low
+ 255.000001n V_hig
+ 255.100000n V_hig
+ 255.100001n V_hig
+ 255.200000n V_hig
+ 255.200001n V_hig
+ 255.300000n V_hig
+ 255.300001n V_hig
+ 255.400000n V_hig
+ 255.400001n V_hig
+ 255.500000n V_hig
+ 255.500001n V_hig
+ 255.600000n V_hig
+ 255.600001n V_hig
+ 255.700000n V_hig
+ 255.700001n V_hig
+ 255.800000n V_hig
+ 255.800001n V_hig
+ 255.900000n V_hig
+ 255.900001n V_hig
+ 256.000000n V_hig
+ 256.000001n V_hig
+ 256.100000n V_hig
+ 256.100001n V_hig
+ 256.200000n V_hig
+ 256.200001n V_hig
+ 256.300000n V_hig
+ 256.300001n V_hig
+ 256.400000n V_hig
+ 256.400001n V_hig
+ 256.500000n V_hig
+ 256.500001n V_hig
+ 256.600000n V_hig
+ 256.600001n V_hig
+ 256.700000n V_hig
+ 256.700001n V_hig
+ 256.800000n V_hig
+ 256.800001n V_hig
+ 256.900000n V_hig
+ 256.900001n V_hig
+ 257.000000n V_hig
+ 257.000001n V_hig
+ 257.100000n V_hig
+ 257.100001n V_hig
+ 257.200000n V_hig
+ 257.200001n V_hig
+ 257.300000n V_hig
+ 257.300001n V_hig
+ 257.400000n V_hig
+ 257.400001n V_hig
+ 257.500000n V_hig
+ 257.500001n V_hig
+ 257.600000n V_hig
+ 257.600001n V_hig
+ 257.700000n V_hig
+ 257.700001n V_hig
+ 257.800000n V_hig
+ 257.800001n V_hig
+ 257.900000n V_hig
+ 257.900001n V_hig
+ 258.000000n V_hig
+ 258.000001n V_hig
+ 258.100000n V_hig
+ 258.100001n V_hig
+ 258.200000n V_hig
+ 258.200001n V_hig
+ 258.300000n V_hig
+ 258.300001n V_hig
+ 258.400000n V_hig
+ 258.400001n V_hig
+ 258.500000n V_hig
+ 258.500001n V_hig
+ 258.600000n V_hig
+ 258.600001n V_hig
+ 258.700000n V_hig
+ 258.700001n V_hig
+ 258.800000n V_hig
+ 258.800001n V_hig
+ 258.900000n V_hig
+ 258.900001n V_hig
+ 259.000000n V_hig
+ 259.000001n V_low
+ 259.100000n V_low
+ 259.100001n V_low
+ 259.200000n V_low
+ 259.200001n V_low
+ 259.300000n V_low
+ 259.300001n V_low
+ 259.400000n V_low
+ 259.400001n V_low
+ 259.500000n V_low
+ 259.500001n V_low
+ 259.600000n V_low
+ 259.600001n V_low
+ 259.700000n V_low
+ 259.700001n V_low
+ 259.800000n V_low
+ 259.800001n V_low
+ 259.900000n V_low
+ 259.900001n V_low
+ 260.000000n V_low
+ 260.000001n V_hig
+ 260.100000n V_hig
+ 260.100001n V_hig
+ 260.200000n V_hig
+ 260.200001n V_hig
+ 260.300000n V_hig
+ 260.300001n V_hig
+ 260.400000n V_hig
+ 260.400001n V_hig
+ 260.500000n V_hig
+ 260.500001n V_hig
+ 260.600000n V_hig
+ 260.600001n V_hig
+ 260.700000n V_hig
+ 260.700001n V_hig
+ 260.800000n V_hig
+ 260.800001n V_hig
+ 260.900000n V_hig
+ 260.900001n V_hig
+ 261.000000n V_hig
+ 261.000001n V_hig
+ 261.100000n V_hig
+ 261.100001n V_hig
+ 261.200000n V_hig
+ 261.200001n V_hig
+ 261.300000n V_hig
+ 261.300001n V_hig
+ 261.400000n V_hig
+ 261.400001n V_hig
+ 261.500000n V_hig
+ 261.500001n V_hig
+ 261.600000n V_hig
+ 261.600001n V_hig
+ 261.700000n V_hig
+ 261.700001n V_hig
+ 261.800000n V_hig
+ 261.800001n V_hig
+ 261.900000n V_hig
+ 261.900001n V_hig
+ 262.000000n V_hig
+ 262.000001n V_hig
+ 262.100000n V_hig
+ 262.100001n V_hig
+ 262.200000n V_hig
+ 262.200001n V_hig
+ 262.300000n V_hig
+ 262.300001n V_hig
+ 262.400000n V_hig
+ 262.400001n V_hig
+ 262.500000n V_hig
+ 262.500001n V_hig
+ 262.600000n V_hig
+ 262.600001n V_hig
+ 262.700000n V_hig
+ 262.700001n V_hig
+ 262.800000n V_hig
+ 262.800001n V_hig
+ 262.900000n V_hig
+ 262.900001n V_hig
+ 263.000000n V_hig
+ 263.000001n V_low
+ 263.100000n V_low
+ 263.100001n V_low
+ 263.200000n V_low
+ 263.200001n V_low
+ 263.300000n V_low
+ 263.300001n V_low
+ 263.400000n V_low
+ 263.400001n V_low
+ 263.500000n V_low
+ 263.500001n V_low
+ 263.600000n V_low
+ 263.600001n V_low
+ 263.700000n V_low
+ 263.700001n V_low
+ 263.800000n V_low
+ 263.800001n V_low
+ 263.900000n V_low
+ 263.900001n V_low
+ 264.000000n V_low
+ 264.000001n V_hig
+ 264.100000n V_hig
+ 264.100001n V_hig
+ 264.200000n V_hig
+ 264.200001n V_hig
+ 264.300000n V_hig
+ 264.300001n V_hig
+ 264.400000n V_hig
+ 264.400001n V_hig
+ 264.500000n V_hig
+ 264.500001n V_hig
+ 264.600000n V_hig
+ 264.600001n V_hig
+ 264.700000n V_hig
+ 264.700001n V_hig
+ 264.800000n V_hig
+ 264.800001n V_hig
+ 264.900000n V_hig
+ 264.900001n V_hig
+ 265.000000n V_hig
+ 265.000001n V_hig
+ 265.100000n V_hig
+ 265.100001n V_hig
+ 265.200000n V_hig
+ 265.200001n V_hig
+ 265.300000n V_hig
+ 265.300001n V_hig
+ 265.400000n V_hig
+ 265.400001n V_hig
+ 265.500000n V_hig
+ 265.500001n V_hig
+ 265.600000n V_hig
+ 265.600001n V_hig
+ 265.700000n V_hig
+ 265.700001n V_hig
+ 265.800000n V_hig
+ 265.800001n V_hig
+ 265.900000n V_hig
+ 265.900001n V_hig
+ 266.000000n V_hig
+ 266.000001n V_low
+ 266.100000n V_low
+ 266.100001n V_low
+ 266.200000n V_low
+ 266.200001n V_low
+ 266.300000n V_low
+ 266.300001n V_low
+ 266.400000n V_low
+ 266.400001n V_low
+ 266.500000n V_low
+ 266.500001n V_low
+ 266.600000n V_low
+ 266.600001n V_low
+ 266.700000n V_low
+ 266.700001n V_low
+ 266.800000n V_low
+ 266.800001n V_low
+ 266.900000n V_low
+ 266.900001n V_low
+ 267.000000n V_low
+ 267.000001n V_low
+ 267.100000n V_low
+ 267.100001n V_low
+ 267.200000n V_low
+ 267.200001n V_low
+ 267.300000n V_low
+ 267.300001n V_low
+ 267.400000n V_low
+ 267.400001n V_low
+ 267.500000n V_low
+ 267.500001n V_low
+ 267.600000n V_low
+ 267.600001n V_low
+ 267.700000n V_low
+ 267.700001n V_low
+ 267.800000n V_low
+ 267.800001n V_low
+ 267.900000n V_low
+ 267.900001n V_low
+ 268.000000n V_low
+ 268.000001n V_low
+ 268.100000n V_low
+ 268.100001n V_low
+ 268.200000n V_low
+ 268.200001n V_low
+ 268.300000n V_low
+ 268.300001n V_low
+ 268.400000n V_low
+ 268.400001n V_low
+ 268.500000n V_low
+ 268.500001n V_low
+ 268.600000n V_low
+ 268.600001n V_low
+ 268.700000n V_low
+ 268.700001n V_low
+ 268.800000n V_low
+ 268.800001n V_low
+ 268.900000n V_low
+ 268.900001n V_low
+ 269.000000n V_low
+ 269.000001n V_low
+ 269.100000n V_low
+ 269.100001n V_low
+ 269.200000n V_low
+ 269.200001n V_low
+ 269.300000n V_low
+ 269.300001n V_low
+ 269.400000n V_low
+ 269.400001n V_low
+ 269.500000n V_low
+ 269.500001n V_low
+ 269.600000n V_low
+ 269.600001n V_low
+ 269.700000n V_low
+ 269.700001n V_low
+ 269.800000n V_low
+ 269.800001n V_low
+ 269.900000n V_low
+ 269.900001n V_low
+ 270.000000n V_low
+ 270.000001n V_hig
+ 270.100000n V_hig
+ 270.100001n V_hig
+ 270.200000n V_hig
+ 270.200001n V_hig
+ 270.300000n V_hig
+ 270.300001n V_hig
+ 270.400000n V_hig
+ 270.400001n V_hig
+ 270.500000n V_hig
+ 270.500001n V_hig
+ 270.600000n V_hig
+ 270.600001n V_hig
+ 270.700000n V_hig
+ 270.700001n V_hig
+ 270.800000n V_hig
+ 270.800001n V_hig
+ 270.900000n V_hig
+ 270.900001n V_hig
+ 271.000000n V_hig
+ 271.000001n V_hig
+ 271.100000n V_hig
+ 271.100001n V_hig
+ 271.200000n V_hig
+ 271.200001n V_hig
+ 271.300000n V_hig
+ 271.300001n V_hig
+ 271.400000n V_hig
+ 271.400001n V_hig
+ 271.500000n V_hig
+ 271.500001n V_hig
+ 271.600000n V_hig
+ 271.600001n V_hig
+ 271.700000n V_hig
+ 271.700001n V_hig
+ 271.800000n V_hig
+ 271.800001n V_hig
+ 271.900000n V_hig
+ 271.900001n V_hig
+ 272.000000n V_hig
+ 272.000001n V_hig
+ 272.100000n V_hig
+ 272.100001n V_hig
+ 272.200000n V_hig
+ 272.200001n V_hig
+ 272.300000n V_hig
+ 272.300001n V_hig
+ 272.400000n V_hig
+ 272.400001n V_hig
+ 272.500000n V_hig
+ 272.500001n V_hig
+ 272.600000n V_hig
+ 272.600001n V_hig
+ 272.700000n V_hig
+ 272.700001n V_hig
+ 272.800000n V_hig
+ 272.800001n V_hig
+ 272.900000n V_hig
+ 272.900001n V_hig
+ 273.000000n V_hig
+ 273.000001n V_hig
+ 273.100000n V_hig
+ 273.100001n V_hig
+ 273.200000n V_hig
+ 273.200001n V_hig
+ 273.300000n V_hig
+ 273.300001n V_hig
+ 273.400000n V_hig
+ 273.400001n V_hig
+ 273.500000n V_hig
+ 273.500001n V_hig
+ 273.600000n V_hig
+ 273.600001n V_hig
+ 273.700000n V_hig
+ 273.700001n V_hig
+ 273.800000n V_hig
+ 273.800001n V_hig
+ 273.900000n V_hig
+ 273.900001n V_hig
+ 274.000000n V_hig
+ 274.000001n V_low
+ 274.100000n V_low
+ 274.100001n V_low
+ 274.200000n V_low
+ 274.200001n V_low
+ 274.300000n V_low
+ 274.300001n V_low
+ 274.400000n V_low
+ 274.400001n V_low
+ 274.500000n V_low
+ 274.500001n V_low
+ 274.600000n V_low
+ 274.600001n V_low
+ 274.700000n V_low
+ 274.700001n V_low
+ 274.800000n V_low
+ 274.800001n V_low
+ 274.900000n V_low
+ 274.900001n V_low
+ 275.000000n V_low
+ 275.000001n V_low
+ 275.100000n V_low
+ 275.100001n V_low
+ 275.200000n V_low
+ 275.200001n V_low
+ 275.300000n V_low
+ 275.300001n V_low
+ 275.400000n V_low
+ 275.400001n V_low
+ 275.500000n V_low
+ 275.500001n V_low
+ 275.600000n V_low
+ 275.600001n V_low
+ 275.700000n V_low
+ 275.700001n V_low
+ 275.800000n V_low
+ 275.800001n V_low
+ 275.900000n V_low
+ 275.900001n V_low
+ 276.000000n V_low
+ 276.000001n V_hig
+ 276.100000n V_hig
+ 276.100001n V_hig
+ 276.200000n V_hig
+ 276.200001n V_hig
+ 276.300000n V_hig
+ 276.300001n V_hig
+ 276.400000n V_hig
+ 276.400001n V_hig
+ 276.500000n V_hig
+ 276.500001n V_hig
+ 276.600000n V_hig
+ 276.600001n V_hig
+ 276.700000n V_hig
+ 276.700001n V_hig
+ 276.800000n V_hig
+ 276.800001n V_hig
+ 276.900000n V_hig
+ 276.900001n V_hig
+ 277.000000n V_hig
+ 277.000001n V_low
+ 277.100000n V_low
+ 277.100001n V_low
+ 277.200000n V_low
+ 277.200001n V_low
+ 277.300000n V_low
+ 277.300001n V_low
+ 277.400000n V_low
+ 277.400001n V_low
+ 277.500000n V_low
+ 277.500001n V_low
+ 277.600000n V_low
+ 277.600001n V_low
+ 277.700000n V_low
+ 277.700001n V_low
+ 277.800000n V_low
+ 277.800001n V_low
+ 277.900000n V_low
+ 277.900001n V_low
+ 278.000000n V_low
+ 278.000001n V_low
+ 278.100000n V_low
+ 278.100001n V_low
+ 278.200000n V_low
+ 278.200001n V_low
+ 278.300000n V_low
+ 278.300001n V_low
+ 278.400000n V_low
+ 278.400001n V_low
+ 278.500000n V_low
+ 278.500001n V_low
+ 278.600000n V_low
+ 278.600001n V_low
+ 278.700000n V_low
+ 278.700001n V_low
+ 278.800000n V_low
+ 278.800001n V_low
+ 278.900000n V_low
+ 278.900001n V_low
+ 279.000000n V_low
+ 279.000001n V_hig
+ 279.100000n V_hig
+ 279.100001n V_hig
+ 279.200000n V_hig
+ 279.200001n V_hig
+ 279.300000n V_hig
+ 279.300001n V_hig
+ 279.400000n V_hig
+ 279.400001n V_hig
+ 279.500000n V_hig
+ 279.500001n V_hig
+ 279.600000n V_hig
+ 279.600001n V_hig
+ 279.700000n V_hig
+ 279.700001n V_hig
+ 279.800000n V_hig
+ 279.800001n V_hig
+ 279.900000n V_hig
+ 279.900001n V_hig
+ 280.000000n V_hig
+ 280.000001n V_hig
+ 280.100000n V_hig
+ 280.100001n V_hig
+ 280.200000n V_hig
+ 280.200001n V_hig
+ 280.300000n V_hig
+ 280.300001n V_hig
+ 280.400000n V_hig
+ 280.400001n V_hig
+ 280.500000n V_hig
+ 280.500001n V_hig
+ 280.600000n V_hig
+ 280.600001n V_hig
+ 280.700000n V_hig
+ 280.700001n V_hig
+ 280.800000n V_hig
+ 280.800001n V_hig
+ 280.900000n V_hig
+ 280.900001n V_hig
+ 281.000000n V_hig
+ 281.000001n V_low
+ 281.100000n V_low
+ 281.100001n V_low
+ 281.200000n V_low
+ 281.200001n V_low
+ 281.300000n V_low
+ 281.300001n V_low
+ 281.400000n V_low
+ 281.400001n V_low
+ 281.500000n V_low
+ 281.500001n V_low
+ 281.600000n V_low
+ 281.600001n V_low
+ 281.700000n V_low
+ 281.700001n V_low
+ 281.800000n V_low
+ 281.800001n V_low
+ 281.900000n V_low
+ 281.900001n V_low
+ 282.000000n V_low
+ 282.000001n V_hig
+ 282.100000n V_hig
+ 282.100001n V_hig
+ 282.200000n V_hig
+ 282.200001n V_hig
+ 282.300000n V_hig
+ 282.300001n V_hig
+ 282.400000n V_hig
+ 282.400001n V_hig
+ 282.500000n V_hig
+ 282.500001n V_hig
+ 282.600000n V_hig
+ 282.600001n V_hig
+ 282.700000n V_hig
+ 282.700001n V_hig
+ 282.800000n V_hig
+ 282.800001n V_hig
+ 282.900000n V_hig
+ 282.900001n V_hig
+ 283.000000n V_hig
+ 283.000001n V_hig
+ 283.100000n V_hig
+ 283.100001n V_hig
+ 283.200000n V_hig
+ 283.200001n V_hig
+ 283.300000n V_hig
+ 283.300001n V_hig
+ 283.400000n V_hig
+ 283.400001n V_hig
+ 283.500000n V_hig
+ 283.500001n V_hig
+ 283.600000n V_hig
+ 283.600001n V_hig
+ 283.700000n V_hig
+ 283.700001n V_hig
+ 283.800000n V_hig
+ 283.800001n V_hig
+ 283.900000n V_hig
+ 283.900001n V_hig
+ 284.000000n V_hig
+ 284.000001n V_hig
+ 284.100000n V_hig
+ 284.100001n V_hig
+ 284.200000n V_hig
+ 284.200001n V_hig
+ 284.300000n V_hig
+ 284.300001n V_hig
+ 284.400000n V_hig
+ 284.400001n V_hig
+ 284.500000n V_hig
+ 284.500001n V_hig
+ 284.600000n V_hig
+ 284.600001n V_hig
+ 284.700000n V_hig
+ 284.700001n V_hig
+ 284.800000n V_hig
+ 284.800001n V_hig
+ 284.900000n V_hig
+ 284.900001n V_hig
+ 285.000000n V_hig
+ 285.000001n V_hig
+ 285.100000n V_hig
+ 285.100001n V_hig
+ 285.200000n V_hig
+ 285.200001n V_hig
+ 285.300000n V_hig
+ 285.300001n V_hig
+ 285.400000n V_hig
+ 285.400001n V_hig
+ 285.500000n V_hig
+ 285.500001n V_hig
+ 285.600000n V_hig
+ 285.600001n V_hig
+ 285.700000n V_hig
+ 285.700001n V_hig
+ 285.800000n V_hig
+ 285.800001n V_hig
+ 285.900000n V_hig
+ 285.900001n V_hig
+ 286.000000n V_hig
+ 286.000001n V_low
+ 286.100000n V_low
+ 286.100001n V_low
+ 286.200000n V_low
+ 286.200001n V_low
+ 286.300000n V_low
+ 286.300001n V_low
+ 286.400000n V_low
+ 286.400001n V_low
+ 286.500000n V_low
+ 286.500001n V_low
+ 286.600000n V_low
+ 286.600001n V_low
+ 286.700000n V_low
+ 286.700001n V_low
+ 286.800000n V_low
+ 286.800001n V_low
+ 286.900000n V_low
+ 286.900001n V_low
+ 287.000000n V_low
+ 287.000001n V_hig
+ 287.100000n V_hig
+ 287.100001n V_hig
+ 287.200000n V_hig
+ 287.200001n V_hig
+ 287.300000n V_hig
+ 287.300001n V_hig
+ 287.400000n V_hig
+ 287.400001n V_hig
+ 287.500000n V_hig
+ 287.500001n V_hig
+ 287.600000n V_hig
+ 287.600001n V_hig
+ 287.700000n V_hig
+ 287.700001n V_hig
+ 287.800000n V_hig
+ 287.800001n V_hig
+ 287.900000n V_hig
+ 287.900001n V_hig
+ 288.000000n V_hig
+ 288.000001n V_hig
+ 288.100000n V_hig
+ 288.100001n V_hig
+ 288.200000n V_hig
+ 288.200001n V_hig
+ 288.300000n V_hig
+ 288.300001n V_hig
+ 288.400000n V_hig
+ 288.400001n V_hig
+ 288.500000n V_hig
+ 288.500001n V_hig
+ 288.600000n V_hig
+ 288.600001n V_hig
+ 288.700000n V_hig
+ 288.700001n V_hig
+ 288.800000n V_hig
+ 288.800001n V_hig
+ 288.900000n V_hig
+ 288.900001n V_hig
+ 289.000000n V_hig
+ 289.000001n V_hig
+ 289.100000n V_hig
+ 289.100001n V_hig
+ 289.200000n V_hig
+ 289.200001n V_hig
+ 289.300000n V_hig
+ 289.300001n V_hig
+ 289.400000n V_hig
+ 289.400001n V_hig
+ 289.500000n V_hig
+ 289.500001n V_hig
+ 289.600000n V_hig
+ 289.600001n V_hig
+ 289.700000n V_hig
+ 289.700001n V_hig
+ 289.800000n V_hig
+ 289.800001n V_hig
+ 289.900000n V_hig
+ 289.900001n V_hig
+ 290.000000n V_hig
+ 290.000001n V_low
+ 290.100000n V_low
+ 290.100001n V_low
+ 290.200000n V_low
+ 290.200001n V_low
+ 290.300000n V_low
+ 290.300001n V_low
+ 290.400000n V_low
+ 290.400001n V_low
+ 290.500000n V_low
+ 290.500001n V_low
+ 290.600000n V_low
+ 290.600001n V_low
+ 290.700000n V_low
+ 290.700001n V_low
+ 290.800000n V_low
+ 290.800001n V_low
+ 290.900000n V_low
+ 290.900001n V_low
+ 291.000000n V_low
+ 291.000001n V_hig
+ 291.100000n V_hig
+ 291.100001n V_hig
+ 291.200000n V_hig
+ 291.200001n V_hig
+ 291.300000n V_hig
+ 291.300001n V_hig
+ 291.400000n V_hig
+ 291.400001n V_hig
+ 291.500000n V_hig
+ 291.500001n V_hig
+ 291.600000n V_hig
+ 291.600001n V_hig
+ 291.700000n V_hig
+ 291.700001n V_hig
+ 291.800000n V_hig
+ 291.800001n V_hig
+ 291.900000n V_hig
+ 291.900001n V_hig
+ 292.000000n V_hig
+ 292.000001n V_hig
+ 292.100000n V_hig
+ 292.100001n V_hig
+ 292.200000n V_hig
+ 292.200001n V_hig
+ 292.300000n V_hig
+ 292.300001n V_hig
+ 292.400000n V_hig
+ 292.400001n V_hig
+ 292.500000n V_hig
+ 292.500001n V_hig
+ 292.600000n V_hig
+ 292.600001n V_hig
+ 292.700000n V_hig
+ 292.700001n V_hig
+ 292.800000n V_hig
+ 292.800001n V_hig
+ 292.900000n V_hig
+ 292.900001n V_hig
+ 293.000000n V_hig
+ 293.000001n V_hig
+ 293.100000n V_hig
+ 293.100001n V_hig
+ 293.200000n V_hig
+ 293.200001n V_hig
+ 293.300000n V_hig
+ 293.300001n V_hig
+ 293.400000n V_hig
+ 293.400001n V_hig
+ 293.500000n V_hig
+ 293.500001n V_hig
+ 293.600000n V_hig
+ 293.600001n V_hig
+ 293.700000n V_hig
+ 293.700001n V_hig
+ 293.800000n V_hig
+ 293.800001n V_hig
+ 293.900000n V_hig
+ 293.900001n V_hig
+ 294.000000n V_hig
+ 294.000001n V_hig
+ 294.100000n V_hig
+ 294.100001n V_hig
+ 294.200000n V_hig
+ 294.200001n V_hig
+ 294.300000n V_hig
+ 294.300001n V_hig
+ 294.400000n V_hig
+ 294.400001n V_hig
+ 294.500000n V_hig
+ 294.500001n V_hig
+ 294.600000n V_hig
+ 294.600001n V_hig
+ 294.700000n V_hig
+ 294.700001n V_hig
+ 294.800000n V_hig
+ 294.800001n V_hig
+ 294.900000n V_hig
+ 294.900001n V_hig
+ 295.000000n V_hig
+ 295.000001n V_low
+ 295.100000n V_low
+ 295.100001n V_low
+ 295.200000n V_low
+ 295.200001n V_low
+ 295.300000n V_low
+ 295.300001n V_low
+ 295.400000n V_low
+ 295.400001n V_low
+ 295.500000n V_low
+ 295.500001n V_low
+ 295.600000n V_low
+ 295.600001n V_low
+ 295.700000n V_low
+ 295.700001n V_low
+ 295.800000n V_low
+ 295.800001n V_low
+ 295.900000n V_low
+ 295.900001n V_low
+ 296.000000n V_low
+ 296.000001n V_low
+ 296.100000n V_low
+ 296.100001n V_low
+ 296.200000n V_low
+ 296.200001n V_low
+ 296.300000n V_low
+ 296.300001n V_low
+ 296.400000n V_low
+ 296.400001n V_low
+ 296.500000n V_low
+ 296.500001n V_low
+ 296.600000n V_low
+ 296.600001n V_low
+ 296.700000n V_low
+ 296.700001n V_low
+ 296.800000n V_low
+ 296.800001n V_low
+ 296.900000n V_low
+ 296.900001n V_low
+ 297.000000n V_low
+ 297.000001n V_low
+ 297.100000n V_low
+ 297.100001n V_low
+ 297.200000n V_low
+ 297.200001n V_low
+ 297.300000n V_low
+ 297.300001n V_low
+ 297.400000n V_low
+ 297.400001n V_low
+ 297.500000n V_low
+ 297.500001n V_low
+ 297.600000n V_low
+ 297.600001n V_low
+ 297.700000n V_low
+ 297.700001n V_low
+ 297.800000n V_low
+ 297.800001n V_low
+ 297.900000n V_low
+ 297.900001n V_low
+ 298.000000n V_low
+ 298.000001n V_low
+ 298.100000n V_low
+ 298.100001n V_low
+ 298.200000n V_low
+ 298.200001n V_low
+ 298.300000n V_low
+ 298.300001n V_low
+ 298.400000n V_low
+ 298.400001n V_low
+ 298.500000n V_low
+ 298.500001n V_low
+ 298.600000n V_low
+ 298.600001n V_low
+ 298.700000n V_low
+ 298.700001n V_low
+ 298.800000n V_low
+ 298.800001n V_low
+ 298.900000n V_low
+ 298.900001n V_low
+ 299.000000n V_low
+ 299.000001n V_low
+ 299.100000n V_low
+ 299.100001n V_low
+ 299.200000n V_low
+ 299.200001n V_low
+ 299.300000n V_low
+ 299.300001n V_low
+ 299.400000n V_low
+ 299.400001n V_low
+ 299.500000n V_low
+ 299.500001n V_low
+ 299.600000n V_low
+ 299.600001n V_low
+ 299.700000n V_low
+ 299.700001n V_low
+ 299.800000n V_low
+ 299.800001n V_low
+ 299.900000n V_low
+ 299.900001n V_low
+ 300.000000n V_low
+ 300.000001n V_hig
+ 300.100000n V_hig
+ 300.100001n V_hig
+ 300.200000n V_hig
+ 300.200001n V_hig
+ 300.300000n V_hig
+ 300.300001n V_hig
+ 300.400000n V_hig
+ 300.400001n V_hig
+ 300.500000n V_hig
+ 300.500001n V_hig
+ 300.600000n V_hig
+ 300.600001n V_hig
+ 300.700000n V_hig
+ 300.700001n V_hig
+ 300.800000n V_hig
+ 300.800001n V_hig
+ 300.900000n V_hig
+ 300.900001n V_hig
+ 301.000000n V_hig
+ 301.000001n V_hig
+ 301.100000n V_hig
+ 301.100001n V_hig
+ 301.200000n V_hig
+ 301.200001n V_hig
+ 301.300000n V_hig
+ 301.300001n V_hig
+ 301.400000n V_hig
+ 301.400001n V_hig
+ 301.500000n V_hig
+ 301.500001n V_hig
+ 301.600000n V_hig
+ 301.600001n V_hig
+ 301.700000n V_hig
+ 301.700001n V_hig
+ 301.800000n V_hig
+ 301.800001n V_hig
+ 301.900000n V_hig
+ 301.900001n V_hig
+ 302.000000n V_hig
+ 302.000001n V_hig
+ 302.100000n V_hig
+ 302.100001n V_hig
+ 302.200000n V_hig
+ 302.200001n V_hig
+ 302.300000n V_hig
+ 302.300001n V_hig
+ 302.400000n V_hig
+ 302.400001n V_hig
+ 302.500000n V_hig
+ 302.500001n V_hig
+ 302.600000n V_hig
+ 302.600001n V_hig
+ 302.700000n V_hig
+ 302.700001n V_hig
+ 302.800000n V_hig
+ 302.800001n V_hig
+ 302.900000n V_hig
+ 302.900001n V_hig
+ 303.000000n V_hig
+ 303.000001n V_low
+ 303.100000n V_low
+ 303.100001n V_low
+ 303.200000n V_low
+ 303.200001n V_low
+ 303.300000n V_low
+ 303.300001n V_low
+ 303.400000n V_low
+ 303.400001n V_low
+ 303.500000n V_low
+ 303.500001n V_low
+ 303.600000n V_low
+ 303.600001n V_low
+ 303.700000n V_low
+ 303.700001n V_low
+ 303.800000n V_low
+ 303.800001n V_low
+ 303.900000n V_low
+ 303.900001n V_low
+ 304.000000n V_low
+ 304.000001n V_hig
+ 304.100000n V_hig
+ 304.100001n V_hig
+ 304.200000n V_hig
+ 304.200001n V_hig
+ 304.300000n V_hig
+ 304.300001n V_hig
+ 304.400000n V_hig
+ 304.400001n V_hig
+ 304.500000n V_hig
+ 304.500001n V_hig
+ 304.600000n V_hig
+ 304.600001n V_hig
+ 304.700000n V_hig
+ 304.700001n V_hig
+ 304.800000n V_hig
+ 304.800001n V_hig
+ 304.900000n V_hig
+ 304.900001n V_hig
+ 305.000000n V_hig
+ 305.000001n V_low
+ 305.100000n V_low
+ 305.100001n V_low
+ 305.200000n V_low
+ 305.200001n V_low
+ 305.300000n V_low
+ 305.300001n V_low
+ 305.400000n V_low
+ 305.400001n V_low
+ 305.500000n V_low
+ 305.500001n V_low
+ 305.600000n V_low
+ 305.600001n V_low
+ 305.700000n V_low
+ 305.700001n V_low
+ 305.800000n V_low
+ 305.800001n V_low
+ 305.900000n V_low
+ 305.900001n V_low
+ 306.000000n V_low
+ 306.000001n V_hig
+ 306.100000n V_hig
+ 306.100001n V_hig
+ 306.200000n V_hig
+ 306.200001n V_hig
+ 306.300000n V_hig
+ 306.300001n V_hig
+ 306.400000n V_hig
+ 306.400001n V_hig
+ 306.500000n V_hig
+ 306.500001n V_hig
+ 306.600000n V_hig
+ 306.600001n V_hig
+ 306.700000n V_hig
+ 306.700001n V_hig
+ 306.800000n V_hig
+ 306.800001n V_hig
+ 306.900000n V_hig
+ 306.900001n V_hig
+ 307.000000n V_hig
+ 307.000001n V_low
+ 307.100000n V_low
+ 307.100001n V_low
+ 307.200000n V_low
+ 307.200001n V_low
+ 307.300000n V_low
+ 307.300001n V_low
+ 307.400000n V_low
+ 307.400001n V_low
+ 307.500000n V_low
+ 307.500001n V_low
+ 307.600000n V_low
+ 307.600001n V_low
+ 307.700000n V_low
+ 307.700001n V_low
+ 307.800000n V_low
+ 307.800001n V_low
+ 307.900000n V_low
+ 307.900001n V_low
+ 308.000000n V_low
+ 308.000001n V_low
+ 308.100000n V_low
+ 308.100001n V_low
+ 308.200000n V_low
+ 308.200001n V_low
+ 308.300000n V_low
+ 308.300001n V_low
+ 308.400000n V_low
+ 308.400001n V_low
+ 308.500000n V_low
+ 308.500001n V_low
+ 308.600000n V_low
+ 308.600001n V_low
+ 308.700000n V_low
+ 308.700001n V_low
+ 308.800000n V_low
+ 308.800001n V_low
+ 308.900000n V_low
+ 308.900001n V_low
+ 309.000000n V_low
+ 309.000001n V_hig
+ 309.100000n V_hig
+ 309.100001n V_hig
+ 309.200000n V_hig
+ 309.200001n V_hig
+ 309.300000n V_hig
+ 309.300001n V_hig
+ 309.400000n V_hig
+ 309.400001n V_hig
+ 309.500000n V_hig
+ 309.500001n V_hig
+ 309.600000n V_hig
+ 309.600001n V_hig
+ 309.700000n V_hig
+ 309.700001n V_hig
+ 309.800000n V_hig
+ 309.800001n V_hig
+ 309.900000n V_hig
+ 309.900001n V_hig
+ 310.000000n V_hig
+ 310.000001n V_low
+ 310.100000n V_low
+ 310.100001n V_low
+ 310.200000n V_low
+ 310.200001n V_low
+ 310.300000n V_low
+ 310.300001n V_low
+ 310.400000n V_low
+ 310.400001n V_low
+ 310.500000n V_low
+ 310.500001n V_low
+ 310.600000n V_low
+ 310.600001n V_low
+ 310.700000n V_low
+ 310.700001n V_low
+ 310.800000n V_low
+ 310.800001n V_low
+ 310.900000n V_low
+ 310.900001n V_low
+ 311.000000n V_low
+ 311.000001n V_hig
+ 311.100000n V_hig
+ 311.100001n V_hig
+ 311.200000n V_hig
+ 311.200001n V_hig
+ 311.300000n V_hig
+ 311.300001n V_hig
+ 311.400000n V_hig
+ 311.400001n V_hig
+ 311.500000n V_hig
+ 311.500001n V_hig
+ 311.600000n V_hig
+ 311.600001n V_hig
+ 311.700000n V_hig
+ 311.700001n V_hig
+ 311.800000n V_hig
+ 311.800001n V_hig
+ 311.900000n V_hig
+ 311.900001n V_hig
+ 312.000000n V_hig
+ 312.000001n V_hig
+ 312.100000n V_hig
+ 312.100001n V_hig
+ 312.200000n V_hig
+ 312.200001n V_hig
+ 312.300000n V_hig
+ 312.300001n V_hig
+ 312.400000n V_hig
+ 312.400001n V_hig
+ 312.500000n V_hig
+ 312.500001n V_hig
+ 312.600000n V_hig
+ 312.600001n V_hig
+ 312.700000n V_hig
+ 312.700001n V_hig
+ 312.800000n V_hig
+ 312.800001n V_hig
+ 312.900000n V_hig
+ 312.900001n V_hig
+ 313.000000n V_hig
+ 313.000001n V_hig
+ 313.100000n V_hig
+ 313.100001n V_hig
+ 313.200000n V_hig
+ 313.200001n V_hig
+ 313.300000n V_hig
+ 313.300001n V_hig
+ 313.400000n V_hig
+ 313.400001n V_hig
+ 313.500000n V_hig
+ 313.500001n V_hig
+ 313.600000n V_hig
+ 313.600001n V_hig
+ 313.700000n V_hig
+ 313.700001n V_hig
+ 313.800000n V_hig
+ 313.800001n V_hig
+ 313.900000n V_hig
+ 313.900001n V_hig
+ 314.000000n V_hig
+ 314.000001n V_hig
+ 314.100000n V_hig
+ 314.100001n V_hig
+ 314.200000n V_hig
+ 314.200001n V_hig
+ 314.300000n V_hig
+ 314.300001n V_hig
+ 314.400000n V_hig
+ 314.400001n V_hig
+ 314.500000n V_hig
+ 314.500001n V_hig
+ 314.600000n V_hig
+ 314.600001n V_hig
+ 314.700000n V_hig
+ 314.700001n V_hig
+ 314.800000n V_hig
+ 314.800001n V_hig
+ 314.900000n V_hig
+ 314.900001n V_hig
+ 315.000000n V_hig
+ 315.000001n V_low
+ 315.100000n V_low
+ 315.100001n V_low
+ 315.200000n V_low
+ 315.200001n V_low
+ 315.300000n V_low
+ 315.300001n V_low
+ 315.400000n V_low
+ 315.400001n V_low
+ 315.500000n V_low
+ 315.500001n V_low
+ 315.600000n V_low
+ 315.600001n V_low
+ 315.700000n V_low
+ 315.700001n V_low
+ 315.800000n V_low
+ 315.800001n V_low
+ 315.900000n V_low
+ 315.900001n V_low
+ 316.000000n V_low
+ 316.000001n V_low
+ 316.100000n V_low
+ 316.100001n V_low
+ 316.200000n V_low
+ 316.200001n V_low
+ 316.300000n V_low
+ 316.300001n V_low
+ 316.400000n V_low
+ 316.400001n V_low
+ 316.500000n V_low
+ 316.500001n V_low
+ 316.600000n V_low
+ 316.600001n V_low
+ 316.700000n V_low
+ 316.700001n V_low
+ 316.800000n V_low
+ 316.800001n V_low
+ 316.900000n V_low
+ 316.900001n V_low
+ 317.000000n V_low
+ 317.000001n V_low
+ 317.100000n V_low
+ 317.100001n V_low
+ 317.200000n V_low
+ 317.200001n V_low
+ 317.300000n V_low
+ 317.300001n V_low
+ 317.400000n V_low
+ 317.400001n V_low
+ 317.500000n V_low
+ 317.500001n V_low
+ 317.600000n V_low
+ 317.600001n V_low
+ 317.700000n V_low
+ 317.700001n V_low
+ 317.800000n V_low
+ 317.800001n V_low
+ 317.900000n V_low
+ 317.900001n V_low
+ 318.000000n V_low
+ 318.000001n V_hig
+ 318.100000n V_hig
+ 318.100001n V_hig
+ 318.200000n V_hig
+ 318.200001n V_hig
+ 318.300000n V_hig
+ 318.300001n V_hig
+ 318.400000n V_hig
+ 318.400001n V_hig
+ 318.500000n V_hig
+ 318.500001n V_hig
+ 318.600000n V_hig
+ 318.600001n V_hig
+ 318.700000n V_hig
+ 318.700001n V_hig
+ 318.800000n V_hig
+ 318.800001n V_hig
+ 318.900000n V_hig
+ 318.900001n V_hig
+ 319.000000n V_hig
+ 319.000001n V_hig
+ 319.100000n V_hig
+ 319.100001n V_hig
+ 319.200000n V_hig
+ 319.200001n V_hig
+ 319.300000n V_hig
+ 319.300001n V_hig
+ 319.400000n V_hig
+ 319.400001n V_hig
+ 319.500000n V_hig
+ 319.500001n V_hig
+ 319.600000n V_hig
+ 319.600001n V_hig
+ 319.700000n V_hig
+ 319.700001n V_hig
+ 319.800000n V_hig
+ 319.800001n V_hig
+ 319.900000n V_hig
+ 319.900001n V_hig
+ 320.000000n V_hig
+ 320.000001n V_hig
+ 320.100000n V_hig
+ 320.100001n V_hig
+ 320.200000n V_hig
+ 320.200001n V_hig
+ 320.300000n V_hig
+ 320.300001n V_hig
+ 320.400000n V_hig
+ 320.400001n V_hig
+ 320.500000n V_hig
+ 320.500001n V_hig
+ 320.600000n V_hig
+ 320.600001n V_hig
+ 320.700000n V_hig
+ 320.700001n V_hig
+ 320.800000n V_hig
+ 320.800001n V_hig
+ 320.900000n V_hig
+ 320.900001n V_hig
+ 321.000000n V_hig
+ 321.000001n V_hig
+ 321.100000n V_hig
+ 321.100001n V_hig
+ 321.200000n V_hig
+ 321.200001n V_hig
+ 321.300000n V_hig
+ 321.300001n V_hig
+ 321.400000n V_hig
+ 321.400001n V_hig
+ 321.500000n V_hig
+ 321.500001n V_hig
+ 321.600000n V_hig
+ 321.600001n V_hig
+ 321.700000n V_hig
+ 321.700001n V_hig
+ 321.800000n V_hig
+ 321.800001n V_hig
+ 321.900000n V_hig
+ 321.900001n V_hig
+ 322.000000n V_hig
+ 322.000001n V_hig
+ 322.100000n V_hig
+ 322.100001n V_hig
+ 322.200000n V_hig
+ 322.200001n V_hig
+ 322.300000n V_hig
+ 322.300001n V_hig
+ 322.400000n V_hig
+ 322.400001n V_hig
+ 322.500000n V_hig
+ 322.500001n V_hig
+ 322.600000n V_hig
+ 322.600001n V_hig
+ 322.700000n V_hig
+ 322.700001n V_hig
+ 322.800000n V_hig
+ 322.800001n V_hig
+ 322.900000n V_hig
+ 322.900001n V_hig
+ 323.000000n V_hig
+ 323.000001n V_low
+ 323.100000n V_low
+ 323.100001n V_low
+ 323.200000n V_low
+ 323.200001n V_low
+ 323.300000n V_low
+ 323.300001n V_low
+ 323.400000n V_low
+ 323.400001n V_low
+ 323.500000n V_low
+ 323.500001n V_low
+ 323.600000n V_low
+ 323.600001n V_low
+ 323.700000n V_low
+ 323.700001n V_low
+ 323.800000n V_low
+ 323.800001n V_low
+ 323.900000n V_low
+ 323.900001n V_low
+ 324.000000n V_low
+ 324.000001n V_hig
+ 324.100000n V_hig
+ 324.100001n V_hig
+ 324.200000n V_hig
+ 324.200001n V_hig
+ 324.300000n V_hig
+ 324.300001n V_hig
+ 324.400000n V_hig
+ 324.400001n V_hig
+ 324.500000n V_hig
+ 324.500001n V_hig
+ 324.600000n V_hig
+ 324.600001n V_hig
+ 324.700000n V_hig
+ 324.700001n V_hig
+ 324.800000n V_hig
+ 324.800001n V_hig
+ 324.900000n V_hig
+ 324.900001n V_hig
+ 325.000000n V_hig
+ 325.000001n V_hig
+ 325.100000n V_hig
+ 325.100001n V_hig
+ 325.200000n V_hig
+ 325.200001n V_hig
+ 325.300000n V_hig
+ 325.300001n V_hig
+ 325.400000n V_hig
+ 325.400001n V_hig
+ 325.500000n V_hig
+ 325.500001n V_hig
+ 325.600000n V_hig
+ 325.600001n V_hig
+ 325.700000n V_hig
+ 325.700001n V_hig
+ 325.800000n V_hig
+ 325.800001n V_hig
+ 325.900000n V_hig
+ 325.900001n V_hig
+ 326.000000n V_hig
+ 326.000001n V_low
+ 326.100000n V_low
+ 326.100001n V_low
+ 326.200000n V_low
+ 326.200001n V_low
+ 326.300000n V_low
+ 326.300001n V_low
+ 326.400000n V_low
+ 326.400001n V_low
+ 326.500000n V_low
+ 326.500001n V_low
+ 326.600000n V_low
+ 326.600001n V_low
+ 326.700000n V_low
+ 326.700001n V_low
+ 326.800000n V_low
+ 326.800001n V_low
+ 326.900000n V_low
+ 326.900001n V_low
+ 327.000000n V_low
+ 327.000001n V_low
+ 327.100000n V_low
+ 327.100001n V_low
+ 327.200000n V_low
+ 327.200001n V_low
+ 327.300000n V_low
+ 327.300001n V_low
+ 327.400000n V_low
+ 327.400001n V_low
+ 327.500000n V_low
+ 327.500001n V_low
+ 327.600000n V_low
+ 327.600001n V_low
+ 327.700000n V_low
+ 327.700001n V_low
+ 327.800000n V_low
+ 327.800001n V_low
+ 327.900000n V_low
+ 327.900001n V_low
+ 328.000000n V_low
+ 328.000001n V_low
+ 328.100000n V_low
+ 328.100001n V_low
+ 328.200000n V_low
+ 328.200001n V_low
+ 328.300000n V_low
+ 328.300001n V_low
+ 328.400000n V_low
+ 328.400001n V_low
+ 328.500000n V_low
+ 328.500001n V_low
+ 328.600000n V_low
+ 328.600001n V_low
+ 328.700000n V_low
+ 328.700001n V_low
+ 328.800000n V_low
+ 328.800001n V_low
+ 328.900000n V_low
+ 328.900001n V_low
+ 329.000000n V_low
+ 329.000001n V_hig
+ 329.100000n V_hig
+ 329.100001n V_hig
+ 329.200000n V_hig
+ 329.200001n V_hig
+ 329.300000n V_hig
+ 329.300001n V_hig
+ 329.400000n V_hig
+ 329.400001n V_hig
+ 329.500000n V_hig
+ 329.500001n V_hig
+ 329.600000n V_hig
+ 329.600001n V_hig
+ 329.700000n V_hig
+ 329.700001n V_hig
+ 329.800000n V_hig
+ 329.800001n V_hig
+ 329.900000n V_hig
+ 329.900001n V_hig
+ 330.000000n V_hig
+ 330.000001n V_low
+ 330.100000n V_low
+ 330.100001n V_low
+ 330.200000n V_low
+ 330.200001n V_low
+ 330.300000n V_low
+ 330.300001n V_low
+ 330.400000n V_low
+ 330.400001n V_low
+ 330.500000n V_low
+ 330.500001n V_low
+ 330.600000n V_low
+ 330.600001n V_low
+ 330.700000n V_low
+ 330.700001n V_low
+ 330.800000n V_low
+ 330.800001n V_low
+ 330.900000n V_low
+ 330.900001n V_low
+ 331.000000n V_low
+ 331.000001n V_low
+ 331.100000n V_low
+ 331.100001n V_low
+ 331.200000n V_low
+ 331.200001n V_low
+ 331.300000n V_low
+ 331.300001n V_low
+ 331.400000n V_low
+ 331.400001n V_low
+ 331.500000n V_low
+ 331.500001n V_low
+ 331.600000n V_low
+ 331.600001n V_low
+ 331.700000n V_low
+ 331.700001n V_low
+ 331.800000n V_low
+ 331.800001n V_low
+ 331.900000n V_low
+ 331.900001n V_low
+ 332.000000n V_low
+ 332.000001n V_hig
+ 332.100000n V_hig
+ 332.100001n V_hig
+ 332.200000n V_hig
+ 332.200001n V_hig
+ 332.300000n V_hig
+ 332.300001n V_hig
+ 332.400000n V_hig
+ 332.400001n V_hig
+ 332.500000n V_hig
+ 332.500001n V_hig
+ 332.600000n V_hig
+ 332.600001n V_hig
+ 332.700000n V_hig
+ 332.700001n V_hig
+ 332.800000n V_hig
+ 332.800001n V_hig
+ 332.900000n V_hig
+ 332.900001n V_hig
+ 333.000000n V_hig
+ 333.000001n V_low
+ 333.100000n V_low
+ 333.100001n V_low
+ 333.200000n V_low
+ 333.200001n V_low
+ 333.300000n V_low
+ 333.300001n V_low
+ 333.400000n V_low
+ 333.400001n V_low
+ 333.500000n V_low
+ 333.500001n V_low
+ 333.600000n V_low
+ 333.600001n V_low
+ 333.700000n V_low
+ 333.700001n V_low
+ 333.800000n V_low
+ 333.800001n V_low
+ 333.900000n V_low
+ 333.900001n V_low
+ 334.000000n V_low
+ 334.000001n V_hig
+ 334.100000n V_hig
+ 334.100001n V_hig
+ 334.200000n V_hig
+ 334.200001n V_hig
+ 334.300000n V_hig
+ 334.300001n V_hig
+ 334.400000n V_hig
+ 334.400001n V_hig
+ 334.500000n V_hig
+ 334.500001n V_hig
+ 334.600000n V_hig
+ 334.600001n V_hig
+ 334.700000n V_hig
+ 334.700001n V_hig
+ 334.800000n V_hig
+ 334.800001n V_hig
+ 334.900000n V_hig
+ 334.900001n V_hig
+ 335.000000n V_hig
+ 335.000001n V_hig
+ 335.100000n V_hig
+ 335.100001n V_hig
+ 335.200000n V_hig
+ 335.200001n V_hig
+ 335.300000n V_hig
+ 335.300001n V_hig
+ 335.400000n V_hig
+ 335.400001n V_hig
+ 335.500000n V_hig
+ 335.500001n V_hig
+ 335.600000n V_hig
+ 335.600001n V_hig
+ 335.700000n V_hig
+ 335.700001n V_hig
+ 335.800000n V_hig
+ 335.800001n V_hig
+ 335.900000n V_hig
+ 335.900001n V_hig
+ 336.000000n V_hig
+ 336.000001n V_low
+ 336.100000n V_low
+ 336.100001n V_low
+ 336.200000n V_low
+ 336.200001n V_low
+ 336.300000n V_low
+ 336.300001n V_low
+ 336.400000n V_low
+ 336.400001n V_low
+ 336.500000n V_low
+ 336.500001n V_low
+ 336.600000n V_low
+ 336.600001n V_low
+ 336.700000n V_low
+ 336.700001n V_low
+ 336.800000n V_low
+ 336.800001n V_low
+ 336.900000n V_low
+ 336.900001n V_low
+ 337.000000n V_low
+ 337.000001n V_low
+ 337.100000n V_low
+ 337.100001n V_low
+ 337.200000n V_low
+ 337.200001n V_low
+ 337.300000n V_low
+ 337.300001n V_low
+ 337.400000n V_low
+ 337.400001n V_low
+ 337.500000n V_low
+ 337.500001n V_low
+ 337.600000n V_low
+ 337.600001n V_low
+ 337.700000n V_low
+ 337.700001n V_low
+ 337.800000n V_low
+ 337.800001n V_low
+ 337.900000n V_low
+ 337.900001n V_low
+ 338.000000n V_low
+ 338.000001n V_hig
+ 338.100000n V_hig
+ 338.100001n V_hig
+ 338.200000n V_hig
+ 338.200001n V_hig
+ 338.300000n V_hig
+ 338.300001n V_hig
+ 338.400000n V_hig
+ 338.400001n V_hig
+ 338.500000n V_hig
+ 338.500001n V_hig
+ 338.600000n V_hig
+ 338.600001n V_hig
+ 338.700000n V_hig
+ 338.700001n V_hig
+ 338.800000n V_hig
+ 338.800001n V_hig
+ 338.900000n V_hig
+ 338.900001n V_hig
+ 339.000000n V_hig
+ 339.000001n V_hig
+ 339.100000n V_hig
+ 339.100001n V_hig
+ 339.200000n V_hig
+ 339.200001n V_hig
+ 339.300000n V_hig
+ 339.300001n V_hig
+ 339.400000n V_hig
+ 339.400001n V_hig
+ 339.500000n V_hig
+ 339.500001n V_hig
+ 339.600000n V_hig
+ 339.600001n V_hig
+ 339.700000n V_hig
+ 339.700001n V_hig
+ 339.800000n V_hig
+ 339.800001n V_hig
+ 339.900000n V_hig
+ 339.900001n V_hig
+ 340.000000n V_hig
+ 340.000001n V_low
+ 340.100000n V_low
+ 340.100001n V_low
+ 340.200000n V_low
+ 340.200001n V_low
+ 340.300000n V_low
+ 340.300001n V_low
+ 340.400000n V_low
+ 340.400001n V_low
+ 340.500000n V_low
+ 340.500001n V_low
+ 340.600000n V_low
+ 340.600001n V_low
+ 340.700000n V_low
+ 340.700001n V_low
+ 340.800000n V_low
+ 340.800001n V_low
+ 340.900000n V_low
+ 340.900001n V_low
+ 341.000000n V_low
+ 341.000001n V_hig
+ 341.100000n V_hig
+ 341.100001n V_hig
+ 341.200000n V_hig
+ 341.200001n V_hig
+ 341.300000n V_hig
+ 341.300001n V_hig
+ 341.400000n V_hig
+ 341.400001n V_hig
+ 341.500000n V_hig
+ 341.500001n V_hig
+ 341.600000n V_hig
+ 341.600001n V_hig
+ 341.700000n V_hig
+ 341.700001n V_hig
+ 341.800000n V_hig
+ 341.800001n V_hig
+ 341.900000n V_hig
+ 341.900001n V_hig
+ 342.000000n V_hig
+ 342.000001n V_low
+ 342.100000n V_low
+ 342.100001n V_low
+ 342.200000n V_low
+ 342.200001n V_low
+ 342.300000n V_low
+ 342.300001n V_low
+ 342.400000n V_low
+ 342.400001n V_low
+ 342.500000n V_low
+ 342.500001n V_low
+ 342.600000n V_low
+ 342.600001n V_low
+ 342.700000n V_low
+ 342.700001n V_low
+ 342.800000n V_low
+ 342.800001n V_low
+ 342.900000n V_low
+ 342.900001n V_low
+ 343.000000n V_low
+ 343.000001n V_low
+ 343.100000n V_low
+ 343.100001n V_low
+ 343.200000n V_low
+ 343.200001n V_low
+ 343.300000n V_low
+ 343.300001n V_low
+ 343.400000n V_low
+ 343.400001n V_low
+ 343.500000n V_low
+ 343.500001n V_low
+ 343.600000n V_low
+ 343.600001n V_low
+ 343.700000n V_low
+ 343.700001n V_low
+ 343.800000n V_low
+ 343.800001n V_low
+ 343.900000n V_low
+ 343.900001n V_low
+ 344.000000n V_low
+ 344.000001n V_low
+ 344.100000n V_low
+ 344.100001n V_low
+ 344.200000n V_low
+ 344.200001n V_low
+ 344.300000n V_low
+ 344.300001n V_low
+ 344.400000n V_low
+ 344.400001n V_low
+ 344.500000n V_low
+ 344.500001n V_low
+ 344.600000n V_low
+ 344.600001n V_low
+ 344.700000n V_low
+ 344.700001n V_low
+ 344.800000n V_low
+ 344.800001n V_low
+ 344.900000n V_low
+ 344.900001n V_low
+ 345.000000n V_low
+ 345.000001n V_hig
+ 345.100000n V_hig
+ 345.100001n V_hig
+ 345.200000n V_hig
+ 345.200001n V_hig
+ 345.300000n V_hig
+ 345.300001n V_hig
+ 345.400000n V_hig
+ 345.400001n V_hig
+ 345.500000n V_hig
+ 345.500001n V_hig
+ 345.600000n V_hig
+ 345.600001n V_hig
+ 345.700000n V_hig
+ 345.700001n V_hig
+ 345.800000n V_hig
+ 345.800001n V_hig
+ 345.900000n V_hig
+ 345.900001n V_hig
+ 346.000000n V_hig
+ 346.000001n V_hig
+ 346.100000n V_hig
+ 346.100001n V_hig
+ 346.200000n V_hig
+ 346.200001n V_hig
+ 346.300000n V_hig
+ 346.300001n V_hig
+ 346.400000n V_hig
+ 346.400001n V_hig
+ 346.500000n V_hig
+ 346.500001n V_hig
+ 346.600000n V_hig
+ 346.600001n V_hig
+ 346.700000n V_hig
+ 346.700001n V_hig
+ 346.800000n V_hig
+ 346.800001n V_hig
+ 346.900000n V_hig
+ 346.900001n V_hig
+ 347.000000n V_hig
+ 347.000001n V_hig
+ 347.100000n V_hig
+ 347.100001n V_hig
+ 347.200000n V_hig
+ 347.200001n V_hig
+ 347.300000n V_hig
+ 347.300001n V_hig
+ 347.400000n V_hig
+ 347.400001n V_hig
+ 347.500000n V_hig
+ 347.500001n V_hig
+ 347.600000n V_hig
+ 347.600001n V_hig
+ 347.700000n V_hig
+ 347.700001n V_hig
+ 347.800000n V_hig
+ 347.800001n V_hig
+ 347.900000n V_hig
+ 347.900001n V_hig
+ 348.000000n V_hig
+ 348.000001n V_low
+ 348.100000n V_low
+ 348.100001n V_low
+ 348.200000n V_low
+ 348.200001n V_low
+ 348.300000n V_low
+ 348.300001n V_low
+ 348.400000n V_low
+ 348.400001n V_low
+ 348.500000n V_low
+ 348.500001n V_low
+ 348.600000n V_low
+ 348.600001n V_low
+ 348.700000n V_low
+ 348.700001n V_low
+ 348.800000n V_low
+ 348.800001n V_low
+ 348.900000n V_low
+ 348.900001n V_low
+ 349.000000n V_low
+ 349.000001n V_hig
+ 349.100000n V_hig
+ 349.100001n V_hig
+ 349.200000n V_hig
+ 349.200001n V_hig
+ 349.300000n V_hig
+ 349.300001n V_hig
+ 349.400000n V_hig
+ 349.400001n V_hig
+ 349.500000n V_hig
+ 349.500001n V_hig
+ 349.600000n V_hig
+ 349.600001n V_hig
+ 349.700000n V_hig
+ 349.700001n V_hig
+ 349.800000n V_hig
+ 349.800001n V_hig
+ 349.900000n V_hig
+ 349.900001n V_hig
+ 350.000000n V_hig
+ 350.000001n V_low
+ 350.100000n V_low
+ 350.100001n V_low
+ 350.200000n V_low
+ 350.200001n V_low
+ 350.300000n V_low
+ 350.300001n V_low
+ 350.400000n V_low
+ 350.400001n V_low
+ 350.500000n V_low
+ 350.500001n V_low
+ 350.600000n V_low
+ 350.600001n V_low
+ 350.700000n V_low
+ 350.700001n V_low
+ 350.800000n V_low
+ 350.800001n V_low
+ 350.900000n V_low
+ 350.900001n V_low
+ 351.000000n V_low
+ 351.000001n V_hig
+ 351.100000n V_hig
+ 351.100001n V_hig
+ 351.200000n V_hig
+ 351.200001n V_hig
+ 351.300000n V_hig
+ 351.300001n V_hig
+ 351.400000n V_hig
+ 351.400001n V_hig
+ 351.500000n V_hig
+ 351.500001n V_hig
+ 351.600000n V_hig
+ 351.600001n V_hig
+ 351.700000n V_hig
+ 351.700001n V_hig
+ 351.800000n V_hig
+ 351.800001n V_hig
+ 351.900000n V_hig
+ 351.900001n V_hig
+ 352.000000n V_hig
+ 352.000001n V_low
+ 352.100000n V_low
+ 352.100001n V_low
+ 352.200000n V_low
+ 352.200001n V_low
+ 352.300000n V_low
+ 352.300001n V_low
+ 352.400000n V_low
+ 352.400001n V_low
+ 352.500000n V_low
+ 352.500001n V_low
+ 352.600000n V_low
+ 352.600001n V_low
+ 352.700000n V_low
+ 352.700001n V_low
+ 352.800000n V_low
+ 352.800001n V_low
+ 352.900000n V_low
+ 352.900001n V_low
+ 353.000000n V_low
+ 353.000001n V_low
+ 353.100000n V_low
+ 353.100001n V_low
+ 353.200000n V_low
+ 353.200001n V_low
+ 353.300000n V_low
+ 353.300001n V_low
+ 353.400000n V_low
+ 353.400001n V_low
+ 353.500000n V_low
+ 353.500001n V_low
+ 353.600000n V_low
+ 353.600001n V_low
+ 353.700000n V_low
+ 353.700001n V_low
+ 353.800000n V_low
+ 353.800001n V_low
+ 353.900000n V_low
+ 353.900001n V_low
+ 354.000000n V_low
+ 354.000001n V_hig
+ 354.100000n V_hig
+ 354.100001n V_hig
+ 354.200000n V_hig
+ 354.200001n V_hig
+ 354.300000n V_hig
+ 354.300001n V_hig
+ 354.400000n V_hig
+ 354.400001n V_hig
+ 354.500000n V_hig
+ 354.500001n V_hig
+ 354.600000n V_hig
+ 354.600001n V_hig
+ 354.700000n V_hig
+ 354.700001n V_hig
+ 354.800000n V_hig
+ 354.800001n V_hig
+ 354.900000n V_hig
+ 354.900001n V_hig
+ 355.000000n V_hig
+ 355.000001n V_low
+ 355.100000n V_low
+ 355.100001n V_low
+ 355.200000n V_low
+ 355.200001n V_low
+ 355.300000n V_low
+ 355.300001n V_low
+ 355.400000n V_low
+ 355.400001n V_low
+ 355.500000n V_low
+ 355.500001n V_low
+ 355.600000n V_low
+ 355.600001n V_low
+ 355.700000n V_low
+ 355.700001n V_low
+ 355.800000n V_low
+ 355.800001n V_low
+ 355.900000n V_low
+ 355.900001n V_low
+ 356.000000n V_low
+ 356.000001n V_hig
+ 356.100000n V_hig
+ 356.100001n V_hig
+ 356.200000n V_hig
+ 356.200001n V_hig
+ 356.300000n V_hig
+ 356.300001n V_hig
+ 356.400000n V_hig
+ 356.400001n V_hig
+ 356.500000n V_hig
+ 356.500001n V_hig
+ 356.600000n V_hig
+ 356.600001n V_hig
+ 356.700000n V_hig
+ 356.700001n V_hig
+ 356.800000n V_hig
+ 356.800001n V_hig
+ 356.900000n V_hig
+ 356.900001n V_hig
+ 357.000000n V_hig
+ 357.000001n V_hig
+ 357.100000n V_hig
+ 357.100001n V_hig
+ 357.200000n V_hig
+ 357.200001n V_hig
+ 357.300000n V_hig
+ 357.300001n V_hig
+ 357.400000n V_hig
+ 357.400001n V_hig
+ 357.500000n V_hig
+ 357.500001n V_hig
+ 357.600000n V_hig
+ 357.600001n V_hig
+ 357.700000n V_hig
+ 357.700001n V_hig
+ 357.800000n V_hig
+ 357.800001n V_hig
+ 357.900000n V_hig
+ 357.900001n V_hig
+ 358.000000n V_hig
+ 358.000001n V_low
+ 358.100000n V_low
+ 358.100001n V_low
+ 358.200000n V_low
+ 358.200001n V_low
+ 358.300000n V_low
+ 358.300001n V_low
+ 358.400000n V_low
+ 358.400001n V_low
+ 358.500000n V_low
+ 358.500001n V_low
+ 358.600000n V_low
+ 358.600001n V_low
+ 358.700000n V_low
+ 358.700001n V_low
+ 358.800000n V_low
+ 358.800001n V_low
+ 358.900000n V_low
+ 358.900001n V_low
+ 359.000000n V_low
+ 359.000001n V_low
+ 359.100000n V_low
+ 359.100001n V_low
+ 359.200000n V_low
+ 359.200001n V_low
+ 359.300000n V_low
+ 359.300001n V_low
+ 359.400000n V_low
+ 359.400001n V_low
+ 359.500000n V_low
+ 359.500001n V_low
+ 359.600000n V_low
+ 359.600001n V_low
+ 359.700000n V_low
+ 359.700001n V_low
+ 359.800000n V_low
+ 359.800001n V_low
+ 359.900000n V_low
+ 359.900001n V_low
+ 360.000000n V_low
+ 360.000001n V_hig
+ 360.100000n V_hig
+ 360.100001n V_hig
+ 360.200000n V_hig
+ 360.200001n V_hig
+ 360.300000n V_hig
+ 360.300001n V_hig
+ 360.400000n V_hig
+ 360.400001n V_hig
+ 360.500000n V_hig
+ 360.500001n V_hig
+ 360.600000n V_hig
+ 360.600001n V_hig
+ 360.700000n V_hig
+ 360.700001n V_hig
+ 360.800000n V_hig
+ 360.800001n V_hig
+ 360.900000n V_hig
+ 360.900001n V_hig
+ 361.000000n V_hig
+ 361.000001n V_low
+ 361.100000n V_low
+ 361.100001n V_low
+ 361.200000n V_low
+ 361.200001n V_low
+ 361.300000n V_low
+ 361.300001n V_low
+ 361.400000n V_low
+ 361.400001n V_low
+ 361.500000n V_low
+ 361.500001n V_low
+ 361.600000n V_low
+ 361.600001n V_low
+ 361.700000n V_low
+ 361.700001n V_low
+ 361.800000n V_low
+ 361.800001n V_low
+ 361.900000n V_low
+ 361.900001n V_low
+ 362.000000n V_low
+ 362.000001n V_hig
+ 362.100000n V_hig
+ 362.100001n V_hig
+ 362.200000n V_hig
+ 362.200001n V_hig
+ 362.300000n V_hig
+ 362.300001n V_hig
+ 362.400000n V_hig
+ 362.400001n V_hig
+ 362.500000n V_hig
+ 362.500001n V_hig
+ 362.600000n V_hig
+ 362.600001n V_hig
+ 362.700000n V_hig
+ 362.700001n V_hig
+ 362.800000n V_hig
+ 362.800001n V_hig
+ 362.900000n V_hig
+ 362.900001n V_hig
+ 363.000000n V_hig
+ 363.000001n V_hig
+ 363.100000n V_hig
+ 363.100001n V_hig
+ 363.200000n V_hig
+ 363.200001n V_hig
+ 363.300000n V_hig
+ 363.300001n V_hig
+ 363.400000n V_hig
+ 363.400001n V_hig
+ 363.500000n V_hig
+ 363.500001n V_hig
+ 363.600000n V_hig
+ 363.600001n V_hig
+ 363.700000n V_hig
+ 363.700001n V_hig
+ 363.800000n V_hig
+ 363.800001n V_hig
+ 363.900000n V_hig
+ 363.900001n V_hig
+ 364.000000n V_hig
+ 364.000001n V_low
+ 364.100000n V_low
+ 364.100001n V_low
+ 364.200000n V_low
+ 364.200001n V_low
+ 364.300000n V_low
+ 364.300001n V_low
+ 364.400000n V_low
+ 364.400001n V_low
+ 364.500000n V_low
+ 364.500001n V_low
+ 364.600000n V_low
+ 364.600001n V_low
+ 364.700000n V_low
+ 364.700001n V_low
+ 364.800000n V_low
+ 364.800001n V_low
+ 364.900000n V_low
+ 364.900001n V_low
+ 365.000000n V_low
+ 365.000001n V_hig
+ 365.100000n V_hig
+ 365.100001n V_hig
+ 365.200000n V_hig
+ 365.200001n V_hig
+ 365.300000n V_hig
+ 365.300001n V_hig
+ 365.400000n V_hig
+ 365.400001n V_hig
+ 365.500000n V_hig
+ 365.500001n V_hig
+ 365.600000n V_hig
+ 365.600001n V_hig
+ 365.700000n V_hig
+ 365.700001n V_hig
+ 365.800000n V_hig
+ 365.800001n V_hig
+ 365.900000n V_hig
+ 365.900001n V_hig
+ 366.000000n V_hig
+ 366.000001n V_hig
+ 366.100000n V_hig
+ 366.100001n V_hig
+ 366.200000n V_hig
+ 366.200001n V_hig
+ 366.300000n V_hig
+ 366.300001n V_hig
+ 366.400000n V_hig
+ 366.400001n V_hig
+ 366.500000n V_hig
+ 366.500001n V_hig
+ 366.600000n V_hig
+ 366.600001n V_hig
+ 366.700000n V_hig
+ 366.700001n V_hig
+ 366.800000n V_hig
+ 366.800001n V_hig
+ 366.900000n V_hig
+ 366.900001n V_hig
+ 367.000000n V_hig
+ 367.000001n V_hig
+ 367.100000n V_hig
+ 367.100001n V_hig
+ 367.200000n V_hig
+ 367.200001n V_hig
+ 367.300000n V_hig
+ 367.300001n V_hig
+ 367.400000n V_hig
+ 367.400001n V_hig
+ 367.500000n V_hig
+ 367.500001n V_hig
+ 367.600000n V_hig
+ 367.600001n V_hig
+ 367.700000n V_hig
+ 367.700001n V_hig
+ 367.800000n V_hig
+ 367.800001n V_hig
+ 367.900000n V_hig
+ 367.900001n V_hig
+ 368.000000n V_hig
+ 368.000001n V_low
+ 368.100000n V_low
+ 368.100001n V_low
+ 368.200000n V_low
+ 368.200001n V_low
+ 368.300000n V_low
+ 368.300001n V_low
+ 368.400000n V_low
+ 368.400001n V_low
+ 368.500000n V_low
+ 368.500001n V_low
+ 368.600000n V_low
+ 368.600001n V_low
+ 368.700000n V_low
+ 368.700001n V_low
+ 368.800000n V_low
+ 368.800001n V_low
+ 368.900000n V_low
+ 368.900001n V_low
+ 369.000000n V_low
+ 369.000001n V_low
+ 369.100000n V_low
+ 369.100001n V_low
+ 369.200000n V_low
+ 369.200001n V_low
+ 369.300000n V_low
+ 369.300001n V_low
+ 369.400000n V_low
+ 369.400001n V_low
+ 369.500000n V_low
+ 369.500001n V_low
+ 369.600000n V_low
+ 369.600001n V_low
+ 369.700000n V_low
+ 369.700001n V_low
+ 369.800000n V_low
+ 369.800001n V_low
+ 369.900000n V_low
+ 369.900001n V_low
+ 370.000000n V_low
+ 370.000001n V_hig
+ 370.100000n V_hig
+ 370.100001n V_hig
+ 370.200000n V_hig
+ 370.200001n V_hig
+ 370.300000n V_hig
+ 370.300001n V_hig
+ 370.400000n V_hig
+ 370.400001n V_hig
+ 370.500000n V_hig
+ 370.500001n V_hig
+ 370.600000n V_hig
+ 370.600001n V_hig
+ 370.700000n V_hig
+ 370.700001n V_hig
+ 370.800000n V_hig
+ 370.800001n V_hig
+ 370.900000n V_hig
+ 370.900001n V_hig
+ 371.000000n V_hig
+ 371.000001n V_low
+ 371.100000n V_low
+ 371.100001n V_low
+ 371.200000n V_low
+ 371.200001n V_low
+ 371.300000n V_low
+ 371.300001n V_low
+ 371.400000n V_low
+ 371.400001n V_low
+ 371.500000n V_low
+ 371.500001n V_low
+ 371.600000n V_low
+ 371.600001n V_low
+ 371.700000n V_low
+ 371.700001n V_low
+ 371.800000n V_low
+ 371.800001n V_low
+ 371.900000n V_low
+ 371.900001n V_low
+ 372.000000n V_low
+ 372.000001n V_hig
+ 372.100000n V_hig
+ 372.100001n V_hig
+ 372.200000n V_hig
+ 372.200001n V_hig
+ 372.300000n V_hig
+ 372.300001n V_hig
+ 372.400000n V_hig
+ 372.400001n V_hig
+ 372.500000n V_hig
+ 372.500001n V_hig
+ 372.600000n V_hig
+ 372.600001n V_hig
+ 372.700000n V_hig
+ 372.700001n V_hig
+ 372.800000n V_hig
+ 372.800001n V_hig
+ 372.900000n V_hig
+ 372.900001n V_hig
+ 373.000000n V_hig
+ 373.000001n V_hig
+ 373.100000n V_hig
+ 373.100001n V_hig
+ 373.200000n V_hig
+ 373.200001n V_hig
+ 373.300000n V_hig
+ 373.300001n V_hig
+ 373.400000n V_hig
+ 373.400001n V_hig
+ 373.500000n V_hig
+ 373.500001n V_hig
+ 373.600000n V_hig
+ 373.600001n V_hig
+ 373.700000n V_hig
+ 373.700001n V_hig
+ 373.800000n V_hig
+ 373.800001n V_hig
+ 373.900000n V_hig
+ 373.900001n V_hig
+ 374.000000n V_hig
+ 374.000001n V_hig
+ 374.100000n V_hig
+ 374.100001n V_hig
+ 374.200000n V_hig
+ 374.200001n V_hig
+ 374.300000n V_hig
+ 374.300001n V_hig
+ 374.400000n V_hig
+ 374.400001n V_hig
+ 374.500000n V_hig
+ 374.500001n V_hig
+ 374.600000n V_hig
+ 374.600001n V_hig
+ 374.700000n V_hig
+ 374.700001n V_hig
+ 374.800000n V_hig
+ 374.800001n V_hig
+ 374.900000n V_hig
+ 374.900001n V_hig
+ 375.000000n V_hig
+ 375.000001n V_low
+ 375.100000n V_low
+ 375.100001n V_low
+ 375.200000n V_low
+ 375.200001n V_low
+ 375.300000n V_low
+ 375.300001n V_low
+ 375.400000n V_low
+ 375.400001n V_low
+ 375.500000n V_low
+ 375.500001n V_low
+ 375.600000n V_low
+ 375.600001n V_low
+ 375.700000n V_low
+ 375.700001n V_low
+ 375.800000n V_low
+ 375.800001n V_low
+ 375.900000n V_low
+ 375.900001n V_low
+ 376.000000n V_low
+ 376.000001n V_hig
+ 376.100000n V_hig
+ 376.100001n V_hig
+ 376.200000n V_hig
+ 376.200001n V_hig
+ 376.300000n V_hig
+ 376.300001n V_hig
+ 376.400000n V_hig
+ 376.400001n V_hig
+ 376.500000n V_hig
+ 376.500001n V_hig
+ 376.600000n V_hig
+ 376.600001n V_hig
+ 376.700000n V_hig
+ 376.700001n V_hig
+ 376.800000n V_hig
+ 376.800001n V_hig
+ 376.900000n V_hig
+ 376.900001n V_hig
+ 377.000000n V_hig
+ 377.000001n V_hig
+ 377.100000n V_hig
+ 377.100001n V_hig
+ 377.200000n V_hig
+ 377.200001n V_hig
+ 377.300000n V_hig
+ 377.300001n V_hig
+ 377.400000n V_hig
+ 377.400001n V_hig
+ 377.500000n V_hig
+ 377.500001n V_hig
+ 377.600000n V_hig
+ 377.600001n V_hig
+ 377.700000n V_hig
+ 377.700001n V_hig
+ 377.800000n V_hig
+ 377.800001n V_hig
+ 377.900000n V_hig
+ 377.900001n V_hig
+ 378.000000n V_hig
+ 378.000001n V_hig
+ 378.100000n V_hig
+ 378.100001n V_hig
+ 378.200000n V_hig
+ 378.200001n V_hig
+ 378.300000n V_hig
+ 378.300001n V_hig
+ 378.400000n V_hig
+ 378.400001n V_hig
+ 378.500000n V_hig
+ 378.500001n V_hig
+ 378.600000n V_hig
+ 378.600001n V_hig
+ 378.700000n V_hig
+ 378.700001n V_hig
+ 378.800000n V_hig
+ 378.800001n V_hig
+ 378.900000n V_hig
+ 378.900001n V_hig
+ 379.000000n V_hig
+ 379.000001n V_low
+ 379.100000n V_low
+ 379.100001n V_low
+ 379.200000n V_low
+ 379.200001n V_low
+ 379.300000n V_low
+ 379.300001n V_low
+ 379.400000n V_low
+ 379.400001n V_low
+ 379.500000n V_low
+ 379.500001n V_low
+ 379.600000n V_low
+ 379.600001n V_low
+ 379.700000n V_low
+ 379.700001n V_low
+ 379.800000n V_low
+ 379.800001n V_low
+ 379.900000n V_low
+ 379.900001n V_low
+ 380.000000n V_low
+ 380.000001n V_hig
+ 380.100000n V_hig
+ 380.100001n V_hig
+ 380.200000n V_hig
+ 380.200001n V_hig
+ 380.300000n V_hig
+ 380.300001n V_hig
+ 380.400000n V_hig
+ 380.400001n V_hig
+ 380.500000n V_hig
+ 380.500001n V_hig
+ 380.600000n V_hig
+ 380.600001n V_hig
+ 380.700000n V_hig
+ 380.700001n V_hig
+ 380.800000n V_hig
+ 380.800001n V_hig
+ 380.900000n V_hig
+ 380.900001n V_hig
+ 381.000000n V_hig
+ 381.000001n V_hig
+ 381.100000n V_hig
+ 381.100001n V_hig
+ 381.200000n V_hig
+ 381.200001n V_hig
+ 381.300000n V_hig
+ 381.300001n V_hig
+ 381.400000n V_hig
+ 381.400001n V_hig
+ 381.500000n V_hig
+ 381.500001n V_hig
+ 381.600000n V_hig
+ 381.600001n V_hig
+ 381.700000n V_hig
+ 381.700001n V_hig
+ 381.800000n V_hig
+ 381.800001n V_hig
+ 381.900000n V_hig
+ 381.900001n V_hig
+ 382.000000n V_hig
+ 382.000001n V_hig
+ 382.100000n V_hig
+ 382.100001n V_hig
+ 382.200000n V_hig
+ 382.200001n V_hig
+ 382.300000n V_hig
+ 382.300001n V_hig
+ 382.400000n V_hig
+ 382.400001n V_hig
+ 382.500000n V_hig
+ 382.500001n V_hig
+ 382.600000n V_hig
+ 382.600001n V_hig
+ 382.700000n V_hig
+ 382.700001n V_hig
+ 382.800000n V_hig
+ 382.800001n V_hig
+ 382.900000n V_hig
+ 382.900001n V_hig
+ 383.000000n V_hig
+ 383.000001n V_low
+ 383.100000n V_low
+ 383.100001n V_low
+ 383.200000n V_low
+ 383.200001n V_low
+ 383.300000n V_low
+ 383.300001n V_low
+ 383.400000n V_low
+ 383.400001n V_low
+ 383.500000n V_low
+ 383.500001n V_low
+ 383.600000n V_low
+ 383.600001n V_low
+ 383.700000n V_low
+ 383.700001n V_low
+ 383.800000n V_low
+ 383.800001n V_low
+ 383.900000n V_low
+ 383.900001n V_low
+ 384.000000n V_low
+ 384.000001n V_low
+ 384.100000n V_low
+ 384.100001n V_low
+ 384.200000n V_low
+ 384.200001n V_low
+ 384.300000n V_low
+ 384.300001n V_low
+ 384.400000n V_low
+ 384.400001n V_low
+ 384.500000n V_low
+ 384.500001n V_low
+ 384.600000n V_low
+ 384.600001n V_low
+ 384.700000n V_low
+ 384.700001n V_low
+ 384.800000n V_low
+ 384.800001n V_low
+ 384.900000n V_low
+ 384.900001n V_low
+ 385.000000n V_low
+ 385.000001n V_low
+ 385.100000n V_low
+ 385.100001n V_low
+ 385.200000n V_low
+ 385.200001n V_low
+ 385.300000n V_low
+ 385.300001n V_low
+ 385.400000n V_low
+ 385.400001n V_low
+ 385.500000n V_low
+ 385.500001n V_low
+ 385.600000n V_low
+ 385.600001n V_low
+ 385.700000n V_low
+ 385.700001n V_low
+ 385.800000n V_low
+ 385.800001n V_low
+ 385.900000n V_low
+ 385.900001n V_low
+ 386.000000n V_low
+ 386.000001n V_low
+ 386.100000n V_low
+ 386.100001n V_low
+ 386.200000n V_low
+ 386.200001n V_low
+ 386.300000n V_low
+ 386.300001n V_low
+ 386.400000n V_low
+ 386.400001n V_low
+ 386.500000n V_low
+ 386.500001n V_low
+ 386.600000n V_low
+ 386.600001n V_low
+ 386.700000n V_low
+ 386.700001n V_low
+ 386.800000n V_low
+ 386.800001n V_low
+ 386.900000n V_low
+ 386.900001n V_low
+ 387.000000n V_low
+ 387.000001n V_hig
+ 387.100000n V_hig
+ 387.100001n V_hig
+ 387.200000n V_hig
+ 387.200001n V_hig
+ 387.300000n V_hig
+ 387.300001n V_hig
+ 387.400000n V_hig
+ 387.400001n V_hig
+ 387.500000n V_hig
+ 387.500001n V_hig
+ 387.600000n V_hig
+ 387.600001n V_hig
+ 387.700000n V_hig
+ 387.700001n V_hig
+ 387.800000n V_hig
+ 387.800001n V_hig
+ 387.900000n V_hig
+ 387.900001n V_hig
+ 388.000000n V_hig
+ 388.000001n V_low
+ 388.100000n V_low
+ 388.100001n V_low
+ 388.200000n V_low
+ 388.200001n V_low
+ 388.300000n V_low
+ 388.300001n V_low
+ 388.400000n V_low
+ 388.400001n V_low
+ 388.500000n V_low
+ 388.500001n V_low
+ 388.600000n V_low
+ 388.600001n V_low
+ 388.700000n V_low
+ 388.700001n V_low
+ 388.800000n V_low
+ 388.800001n V_low
+ 388.900000n V_low
+ 388.900001n V_low
+ 389.000000n V_low
+ 389.000001n V_low
+ 389.100000n V_low
+ 389.100001n V_low
+ 389.200000n V_low
+ 389.200001n V_low
+ 389.300000n V_low
+ 389.300001n V_low
+ 389.400000n V_low
+ 389.400001n V_low
+ 389.500000n V_low
+ 389.500001n V_low
+ 389.600000n V_low
+ 389.600001n V_low
+ 389.700000n V_low
+ 389.700001n V_low
+ 389.800000n V_low
+ 389.800001n V_low
+ 389.900000n V_low
+ 389.900001n V_low
+ 390.000000n V_low
+ 390.000001n V_low
+ 390.100000n V_low
+ 390.100001n V_low
+ 390.200000n V_low
+ 390.200001n V_low
+ 390.300000n V_low
+ 390.300001n V_low
+ 390.400000n V_low
+ 390.400001n V_low
+ 390.500000n V_low
+ 390.500001n V_low
+ 390.600000n V_low
+ 390.600001n V_low
+ 390.700000n V_low
+ 390.700001n V_low
+ 390.800000n V_low
+ 390.800001n V_low
+ 390.900000n V_low
+ 390.900001n V_low
+ 391.000000n V_low
+ 391.000001n V_low
+ 391.100000n V_low
+ 391.100001n V_low
+ 391.200000n V_low
+ 391.200001n V_low
+ 391.300000n V_low
+ 391.300001n V_low
+ 391.400000n V_low
+ 391.400001n V_low
+ 391.500000n V_low
+ 391.500001n V_low
+ 391.600000n V_low
+ 391.600001n V_low
+ 391.700000n V_low
+ 391.700001n V_low
+ 391.800000n V_low
+ 391.800001n V_low
+ 391.900000n V_low
+ 391.900001n V_low
+ 392.000000n V_low
+ 392.000001n V_hig
+ 392.100000n V_hig
+ 392.100001n V_hig
+ 392.200000n V_hig
+ 392.200001n V_hig
+ 392.300000n V_hig
+ 392.300001n V_hig
+ 392.400000n V_hig
+ 392.400001n V_hig
+ 392.500000n V_hig
+ 392.500001n V_hig
+ 392.600000n V_hig
+ 392.600001n V_hig
+ 392.700000n V_hig
+ 392.700001n V_hig
+ 392.800000n V_hig
+ 392.800001n V_hig
+ 392.900000n V_hig
+ 392.900001n V_hig
+ 393.000000n V_hig
+ 393.000001n V_low
+ 393.100000n V_low
+ 393.100001n V_low
+ 393.200000n V_low
+ 393.200001n V_low
+ 393.300000n V_low
+ 393.300001n V_low
+ 393.400000n V_low
+ 393.400001n V_low
+ 393.500000n V_low
+ 393.500001n V_low
+ 393.600000n V_low
+ 393.600001n V_low
+ 393.700000n V_low
+ 393.700001n V_low
+ 393.800000n V_low
+ 393.800001n V_low
+ 393.900000n V_low
+ 393.900001n V_low
+ 394.000000n V_low
+ 394.000001n V_hig
+ 394.100000n V_hig
+ 394.100001n V_hig
+ 394.200000n V_hig
+ 394.200001n V_hig
+ 394.300000n V_hig
+ 394.300001n V_hig
+ 394.400000n V_hig
+ 394.400001n V_hig
+ 394.500000n V_hig
+ 394.500001n V_hig
+ 394.600000n V_hig
+ 394.600001n V_hig
+ 394.700000n V_hig
+ 394.700001n V_hig
+ 394.800000n V_hig
+ 394.800001n V_hig
+ 394.900000n V_hig
+ 394.900001n V_hig
+ 395.000000n V_hig
+ 395.000001n V_hig
+ 395.100000n V_hig
+ 395.100001n V_hig
+ 395.200000n V_hig
+ 395.200001n V_hig
+ 395.300000n V_hig
+ 395.300001n V_hig
+ 395.400000n V_hig
+ 395.400001n V_hig
+ 395.500000n V_hig
+ 395.500001n V_hig
+ 395.600000n V_hig
+ 395.600001n V_hig
+ 395.700000n V_hig
+ 395.700001n V_hig
+ 395.800000n V_hig
+ 395.800001n V_hig
+ 395.900000n V_hig
+ 395.900001n V_hig
+ 396.000000n V_hig
+ 396.000001n V_low
+ 396.100000n V_low
+ 396.100001n V_low
+ 396.200000n V_low
+ 396.200001n V_low
+ 396.300000n V_low
+ 396.300001n V_low
+ 396.400000n V_low
+ 396.400001n V_low
+ 396.500000n V_low
+ 396.500001n V_low
+ 396.600000n V_low
+ 396.600001n V_low
+ 396.700000n V_low
+ 396.700001n V_low
+ 396.800000n V_low
+ 396.800001n V_low
+ 396.900000n V_low
+ 396.900001n V_low
+ 397.000000n V_low
+ 397.000001n V_low
+ 397.100000n V_low
+ 397.100001n V_low
+ 397.200000n V_low
+ 397.200001n V_low
+ 397.300000n V_low
+ 397.300001n V_low
+ 397.400000n V_low
+ 397.400001n V_low
+ 397.500000n V_low
+ 397.500001n V_low
+ 397.600000n V_low
+ 397.600001n V_low
+ 397.700000n V_low
+ 397.700001n V_low
+ 397.800000n V_low
+ 397.800001n V_low
+ 397.900000n V_low
+ 397.900001n V_low
+ 398.000000n V_low
+ 398.000001n V_hig
+ 398.100000n V_hig
+ 398.100001n V_hig
+ 398.200000n V_hig
+ 398.200001n V_hig
+ 398.300000n V_hig
+ 398.300001n V_hig
+ 398.400000n V_hig
+ 398.400001n V_hig
+ 398.500000n V_hig
+ 398.500001n V_hig
+ 398.600000n V_hig
+ 398.600001n V_hig
+ 398.700000n V_hig
+ 398.700001n V_hig
+ 398.800000n V_hig
+ 398.800001n V_hig
+ 398.900000n V_hig
+ 398.900001n V_hig
+ 399.000000n V_hig
+ 399.000001n V_low
+ 399.100000n V_low
+ 399.100001n V_low
+ 399.200000n V_low
+ 399.200001n V_low
+ 399.300000n V_low
+ 399.300001n V_low
+ 399.400000n V_low
+ 399.400001n V_low
+ 399.500000n V_low
+ 399.500001n V_low
+ 399.600000n V_low
+ 399.600001n V_low
+ 399.700000n V_low
+ 399.700001n V_low
+ 399.800000n V_low
+ 399.800001n V_low
+ 399.900000n V_low
+ 399.900001n V_low
+ 400.000000n V_low
+ 400.000001n V_hig
+ 400.100000n V_hig
+ 400.100001n V_hig
+ 400.200000n V_hig
+ 400.200001n V_hig
+ 400.300000n V_hig
+ 400.300001n V_hig
+ 400.400000n V_hig
+ 400.400001n V_hig
+ 400.500000n V_hig
+ 400.500001n V_hig
+ 400.600000n V_hig
+ 400.600001n V_hig
+ 400.700000n V_hig
+ 400.700001n V_hig
+ 400.800000n V_hig
+ 400.800001n V_hig
+ 400.900000n V_hig
+ 400.900001n V_hig
+ 401.000000n V_hig
+ 401.000001n V_low
+ 401.100000n V_low
+ 401.100001n V_low
+ 401.200000n V_low
+ 401.200001n V_low
+ 401.300000n V_low
+ 401.300001n V_low
+ 401.400000n V_low
+ 401.400001n V_low
+ 401.500000n V_low
+ 401.500001n V_low
+ 401.600000n V_low
+ 401.600001n V_low
+ 401.700000n V_low
+ 401.700001n V_low
+ 401.800000n V_low
+ 401.800001n V_low
+ 401.900000n V_low
+ 401.900001n V_low
+ 402.000000n V_low
+ 402.000001n V_hig
+ 402.100000n V_hig
+ 402.100001n V_hig
+ 402.200000n V_hig
+ 402.200001n V_hig
+ 402.300000n V_hig
+ 402.300001n V_hig
+ 402.400000n V_hig
+ 402.400001n V_hig
+ 402.500000n V_hig
+ 402.500001n V_hig
+ 402.600000n V_hig
+ 402.600001n V_hig
+ 402.700000n V_hig
+ 402.700001n V_hig
+ 402.800000n V_hig
+ 402.800001n V_hig
+ 402.900000n V_hig
+ 402.900001n V_hig
+ 403.000000n V_hig
+ 403.000001n V_hig
+ 403.100000n V_hig
+ 403.100001n V_hig
+ 403.200000n V_hig
+ 403.200001n V_hig
+ 403.300000n V_hig
+ 403.300001n V_hig
+ 403.400000n V_hig
+ 403.400001n V_hig
+ 403.500000n V_hig
+ 403.500001n V_hig
+ 403.600000n V_hig
+ 403.600001n V_hig
+ 403.700000n V_hig
+ 403.700001n V_hig
+ 403.800000n V_hig
+ 403.800001n V_hig
+ 403.900000n V_hig
+ 403.900001n V_hig
+ 404.000000n V_hig
+ 404.000001n V_hig
+ 404.100000n V_hig
+ 404.100001n V_hig
+ 404.200000n V_hig
+ 404.200001n V_hig
+ 404.300000n V_hig
+ 404.300001n V_hig
+ 404.400000n V_hig
+ 404.400001n V_hig
+ 404.500000n V_hig
+ 404.500001n V_hig
+ 404.600000n V_hig
+ 404.600001n V_hig
+ 404.700000n V_hig
+ 404.700001n V_hig
+ 404.800000n V_hig
+ 404.800001n V_hig
+ 404.900000n V_hig
+ 404.900001n V_hig
+ 405.000000n V_hig
+ 405.000001n V_low
+ 405.100000n V_low
+ 405.100001n V_low
+ 405.200000n V_low
+ 405.200001n V_low
+ 405.300000n V_low
+ 405.300001n V_low
+ 405.400000n V_low
+ 405.400001n V_low
+ 405.500000n V_low
+ 405.500001n V_low
+ 405.600000n V_low
+ 405.600001n V_low
+ 405.700000n V_low
+ 405.700001n V_low
+ 405.800000n V_low
+ 405.800001n V_low
+ 405.900000n V_low
+ 405.900001n V_low
+ 406.000000n V_low
+ 406.000001n V_low
+ 406.100000n V_low
+ 406.100001n V_low
+ 406.200000n V_low
+ 406.200001n V_low
+ 406.300000n V_low
+ 406.300001n V_low
+ 406.400000n V_low
+ 406.400001n V_low
+ 406.500000n V_low
+ 406.500001n V_low
+ 406.600000n V_low
+ 406.600001n V_low
+ 406.700000n V_low
+ 406.700001n V_low
+ 406.800000n V_low
+ 406.800001n V_low
+ 406.900000n V_low
+ 406.900001n V_low
+ 407.000000n V_low
+ 407.000001n V_low
+ 407.100000n V_low
+ 407.100001n V_low
+ 407.200000n V_low
+ 407.200001n V_low
+ 407.300000n V_low
+ 407.300001n V_low
+ 407.400000n V_low
+ 407.400001n V_low
+ 407.500000n V_low
+ 407.500001n V_low
+ 407.600000n V_low
+ 407.600001n V_low
+ 407.700000n V_low
+ 407.700001n V_low
+ 407.800000n V_low
+ 407.800001n V_low
+ 407.900000n V_low
+ 407.900001n V_low
+ 408.000000n V_low
+ 408.000001n V_hig
+ 408.100000n V_hig
+ 408.100001n V_hig
+ 408.200000n V_hig
+ 408.200001n V_hig
+ 408.300000n V_hig
+ 408.300001n V_hig
+ 408.400000n V_hig
+ 408.400001n V_hig
+ 408.500000n V_hig
+ 408.500001n V_hig
+ 408.600000n V_hig
+ 408.600001n V_hig
+ 408.700000n V_hig
+ 408.700001n V_hig
+ 408.800000n V_hig
+ 408.800001n V_hig
+ 408.900000n V_hig
+ 408.900001n V_hig
+ 409.000000n V_hig
+ 409.000001n V_low
+ 409.100000n V_low
+ 409.100001n V_low
+ 409.200000n V_low
+ 409.200001n V_low
+ 409.300000n V_low
+ 409.300001n V_low
+ 409.400000n V_low
+ 409.400001n V_low
+ 409.500000n V_low
+ 409.500001n V_low
+ 409.600000n V_low
+ 409.600001n V_low
+ 409.700000n V_low
+ 409.700001n V_low
+ 409.800000n V_low
+ 409.800001n V_low
+ 409.900000n V_low
+ 409.900001n V_low
+ 410.000000n V_low
+ 410.000001n V_hig
+ 410.100000n V_hig
+ 410.100001n V_hig
+ 410.200000n V_hig
+ 410.200001n V_hig
+ 410.300000n V_hig
+ 410.300001n V_hig
+ 410.400000n V_hig
+ 410.400001n V_hig
+ 410.500000n V_hig
+ 410.500001n V_hig
+ 410.600000n V_hig
+ 410.600001n V_hig
+ 410.700000n V_hig
+ 410.700001n V_hig
+ 410.800000n V_hig
+ 410.800001n V_hig
+ 410.900000n V_hig
+ 410.900001n V_hig
+ 411.000000n V_hig
+ 411.000001n V_low
+ 411.100000n V_low
+ 411.100001n V_low
+ 411.200000n V_low
+ 411.200001n V_low
+ 411.300000n V_low
+ 411.300001n V_low
+ 411.400000n V_low
+ 411.400001n V_low
+ 411.500000n V_low
+ 411.500001n V_low
+ 411.600000n V_low
+ 411.600001n V_low
+ 411.700000n V_low
+ 411.700001n V_low
+ 411.800000n V_low
+ 411.800001n V_low
+ 411.900000n V_low
+ 411.900001n V_low
+ 412.000000n V_low
+ 412.000001n V_low
+ 412.100000n V_low
+ 412.100001n V_low
+ 412.200000n V_low
+ 412.200001n V_low
+ 412.300000n V_low
+ 412.300001n V_low
+ 412.400000n V_low
+ 412.400001n V_low
+ 412.500000n V_low
+ 412.500001n V_low
+ 412.600000n V_low
+ 412.600001n V_low
+ 412.700000n V_low
+ 412.700001n V_low
+ 412.800000n V_low
+ 412.800001n V_low
+ 412.900000n V_low
+ 412.900001n V_low
+ 413.000000n V_low
+ 413.000001n V_low
+ 413.100000n V_low
+ 413.100001n V_low
+ 413.200000n V_low
+ 413.200001n V_low
+ 413.300000n V_low
+ 413.300001n V_low
+ 413.400000n V_low
+ 413.400001n V_low
+ 413.500000n V_low
+ 413.500001n V_low
+ 413.600000n V_low
+ 413.600001n V_low
+ 413.700000n V_low
+ 413.700001n V_low
+ 413.800000n V_low
+ 413.800001n V_low
+ 413.900000n V_low
+ 413.900001n V_low
+ 414.000000n V_low
+ 414.000001n V_hig
+ 414.100000n V_hig
+ 414.100001n V_hig
+ 414.200000n V_hig
+ 414.200001n V_hig
+ 414.300000n V_hig
+ 414.300001n V_hig
+ 414.400000n V_hig
+ 414.400001n V_hig
+ 414.500000n V_hig
+ 414.500001n V_hig
+ 414.600000n V_hig
+ 414.600001n V_hig
+ 414.700000n V_hig
+ 414.700001n V_hig
+ 414.800000n V_hig
+ 414.800001n V_hig
+ 414.900000n V_hig
+ 414.900001n V_hig
+ 415.000000n V_hig
+ 415.000001n V_low
+ 415.100000n V_low
+ 415.100001n V_low
+ 415.200000n V_low
+ 415.200001n V_low
+ 415.300000n V_low
+ 415.300001n V_low
+ 415.400000n V_low
+ 415.400001n V_low
+ 415.500000n V_low
+ 415.500001n V_low
+ 415.600000n V_low
+ 415.600001n V_low
+ 415.700000n V_low
+ 415.700001n V_low
+ 415.800000n V_low
+ 415.800001n V_low
+ 415.900000n V_low
+ 415.900001n V_low
+ 416.000000n V_low
+ 416.000001n V_hig
+ 416.100000n V_hig
+ 416.100001n V_hig
+ 416.200000n V_hig
+ 416.200001n V_hig
+ 416.300000n V_hig
+ 416.300001n V_hig
+ 416.400000n V_hig
+ 416.400001n V_hig
+ 416.500000n V_hig
+ 416.500001n V_hig
+ 416.600000n V_hig
+ 416.600001n V_hig
+ 416.700000n V_hig
+ 416.700001n V_hig
+ 416.800000n V_hig
+ 416.800001n V_hig
+ 416.900000n V_hig
+ 416.900001n V_hig
+ 417.000000n V_hig
+ 417.000001n V_low
+ 417.100000n V_low
+ 417.100001n V_low
+ 417.200000n V_low
+ 417.200001n V_low
+ 417.300000n V_low
+ 417.300001n V_low
+ 417.400000n V_low
+ 417.400001n V_low
+ 417.500000n V_low
+ 417.500001n V_low
+ 417.600000n V_low
+ 417.600001n V_low
+ 417.700000n V_low
+ 417.700001n V_low
+ 417.800000n V_low
+ 417.800001n V_low
+ 417.900000n V_low
+ 417.900001n V_low
+ 418.000000n V_low
+ 418.000001n V_hig
+ 418.100000n V_hig
+ 418.100001n V_hig
+ 418.200000n V_hig
+ 418.200001n V_hig
+ 418.300000n V_hig
+ 418.300001n V_hig
+ 418.400000n V_hig
+ 418.400001n V_hig
+ 418.500000n V_hig
+ 418.500001n V_hig
+ 418.600000n V_hig
+ 418.600001n V_hig
+ 418.700000n V_hig
+ 418.700001n V_hig
+ 418.800000n V_hig
+ 418.800001n V_hig
+ 418.900000n V_hig
+ 418.900001n V_hig
+ 419.000000n V_hig
+ 419.000001n V_hig
+ 419.100000n V_hig
+ 419.100001n V_hig
+ 419.200000n V_hig
+ 419.200001n V_hig
+ 419.300000n V_hig
+ 419.300001n V_hig
+ 419.400000n V_hig
+ 419.400001n V_hig
+ 419.500000n V_hig
+ 419.500001n V_hig
+ 419.600000n V_hig
+ 419.600001n V_hig
+ 419.700000n V_hig
+ 419.700001n V_hig
+ 419.800000n V_hig
+ 419.800001n V_hig
+ 419.900000n V_hig
+ 419.900001n V_hig
+ 420.000000n V_hig
+ 420.000001n V_low
+ 420.100000n V_low
+ 420.100001n V_low
+ 420.200000n V_low
+ 420.200001n V_low
+ 420.300000n V_low
+ 420.300001n V_low
+ 420.400000n V_low
+ 420.400001n V_low
+ 420.500000n V_low
+ 420.500001n V_low
+ 420.600000n V_low
+ 420.600001n V_low
+ 420.700000n V_low
+ 420.700001n V_low
+ 420.800000n V_low
+ 420.800001n V_low
+ 420.900000n V_low
+ 420.900001n V_low
+ 421.000000n V_low
+ 421.000001n V_hig
+ 421.100000n V_hig
+ 421.100001n V_hig
+ 421.200000n V_hig
+ 421.200001n V_hig
+ 421.300000n V_hig
+ 421.300001n V_hig
+ 421.400000n V_hig
+ 421.400001n V_hig
+ 421.500000n V_hig
+ 421.500001n V_hig
+ 421.600000n V_hig
+ 421.600001n V_hig
+ 421.700000n V_hig
+ 421.700001n V_hig
+ 421.800000n V_hig
+ 421.800001n V_hig
+ 421.900000n V_hig
+ 421.900001n V_hig
+ 422.000000n V_hig
+ 422.000001n V_low
+ 422.100000n V_low
+ 422.100001n V_low
+ 422.200000n V_low
+ 422.200001n V_low
+ 422.300000n V_low
+ 422.300001n V_low
+ 422.400000n V_low
+ 422.400001n V_low
+ 422.500000n V_low
+ 422.500001n V_low
+ 422.600000n V_low
+ 422.600001n V_low
+ 422.700000n V_low
+ 422.700001n V_low
+ 422.800000n V_low
+ 422.800001n V_low
+ 422.900000n V_low
+ 422.900001n V_low
+ 423.000000n V_low
+ 423.000001n V_low
+ 423.100000n V_low
+ 423.100001n V_low
+ 423.200000n V_low
+ 423.200001n V_low
+ 423.300000n V_low
+ 423.300001n V_low
+ 423.400000n V_low
+ 423.400001n V_low
+ 423.500000n V_low
+ 423.500001n V_low
+ 423.600000n V_low
+ 423.600001n V_low
+ 423.700000n V_low
+ 423.700001n V_low
+ 423.800000n V_low
+ 423.800001n V_low
+ 423.900000n V_low
+ 423.900001n V_low
+ 424.000000n V_low
+ 424.000001n V_low
+ 424.100000n V_low
+ 424.100001n V_low
+ 424.200000n V_low
+ 424.200001n V_low
+ 424.300000n V_low
+ 424.300001n V_low
+ 424.400000n V_low
+ 424.400001n V_low
+ 424.500000n V_low
+ 424.500001n V_low
+ 424.600000n V_low
+ 424.600001n V_low
+ 424.700000n V_low
+ 424.700001n V_low
+ 424.800000n V_low
+ 424.800001n V_low
+ 424.900000n V_low
+ 424.900001n V_low
+ 425.000000n V_low
+ 425.000001n V_hig
+ 425.100000n V_hig
+ 425.100001n V_hig
+ 425.200000n V_hig
+ 425.200001n V_hig
+ 425.300000n V_hig
+ 425.300001n V_hig
+ 425.400000n V_hig
+ 425.400001n V_hig
+ 425.500000n V_hig
+ 425.500001n V_hig
+ 425.600000n V_hig
+ 425.600001n V_hig
+ 425.700000n V_hig
+ 425.700001n V_hig
+ 425.800000n V_hig
+ 425.800001n V_hig
+ 425.900000n V_hig
+ 425.900001n V_hig
+ 426.000000n V_hig
+ 426.000001n V_hig
+ 426.100000n V_hig
+ 426.100001n V_hig
+ 426.200000n V_hig
+ 426.200001n V_hig
+ 426.300000n V_hig
+ 426.300001n V_hig
+ 426.400000n V_hig
+ 426.400001n V_hig
+ 426.500000n V_hig
+ 426.500001n V_hig
+ 426.600000n V_hig
+ 426.600001n V_hig
+ 426.700000n V_hig
+ 426.700001n V_hig
+ 426.800000n V_hig
+ 426.800001n V_hig
+ 426.900000n V_hig
+ 426.900001n V_hig
+ 427.000000n V_hig
+ 427.000001n V_hig
+ 427.100000n V_hig
+ 427.100001n V_hig
+ 427.200000n V_hig
+ 427.200001n V_hig
+ 427.300000n V_hig
+ 427.300001n V_hig
+ 427.400000n V_hig
+ 427.400001n V_hig
+ 427.500000n V_hig
+ 427.500001n V_hig
+ 427.600000n V_hig
+ 427.600001n V_hig
+ 427.700000n V_hig
+ 427.700001n V_hig
+ 427.800000n V_hig
+ 427.800001n V_hig
+ 427.900000n V_hig
+ 427.900001n V_hig
+ 428.000000n V_hig
+ 428.000001n V_hig
+ 428.100000n V_hig
+ 428.100001n V_hig
+ 428.200000n V_hig
+ 428.200001n V_hig
+ 428.300000n V_hig
+ 428.300001n V_hig
+ 428.400000n V_hig
+ 428.400001n V_hig
+ 428.500000n V_hig
+ 428.500001n V_hig
+ 428.600000n V_hig
+ 428.600001n V_hig
+ 428.700000n V_hig
+ 428.700001n V_hig
+ 428.800000n V_hig
+ 428.800001n V_hig
+ 428.900000n V_hig
+ 428.900001n V_hig
+ 429.000000n V_hig
+ 429.000001n V_hig
+ 429.100000n V_hig
+ 429.100001n V_hig
+ 429.200000n V_hig
+ 429.200001n V_hig
+ 429.300000n V_hig
+ 429.300001n V_hig
+ 429.400000n V_hig
+ 429.400001n V_hig
+ 429.500000n V_hig
+ 429.500001n V_hig
+ 429.600000n V_hig
+ 429.600001n V_hig
+ 429.700000n V_hig
+ 429.700001n V_hig
+ 429.800000n V_hig
+ 429.800001n V_hig
+ 429.900000n V_hig
+ 429.900001n V_hig
+ 430.000000n V_hig
+ 430.000001n V_low
+ 430.100000n V_low
+ 430.100001n V_low
+ 430.200000n V_low
+ 430.200001n V_low
+ 430.300000n V_low
+ 430.300001n V_low
+ 430.400000n V_low
+ 430.400001n V_low
+ 430.500000n V_low
+ 430.500001n V_low
+ 430.600000n V_low
+ 430.600001n V_low
+ 430.700000n V_low
+ 430.700001n V_low
+ 430.800000n V_low
+ 430.800001n V_low
+ 430.900000n V_low
+ 430.900001n V_low
+ 431.000000n V_low
+ 431.000001n V_low
+ 431.100000n V_low
+ 431.100001n V_low
+ 431.200000n V_low
+ 431.200001n V_low
+ 431.300000n V_low
+ 431.300001n V_low
+ 431.400000n V_low
+ 431.400001n V_low
+ 431.500000n V_low
+ 431.500001n V_low
+ 431.600000n V_low
+ 431.600001n V_low
+ 431.700000n V_low
+ 431.700001n V_low
+ 431.800000n V_low
+ 431.800001n V_low
+ 431.900000n V_low
+ 431.900001n V_low
+ 432.000000n V_low
+ 432.000001n V_hig
+ 432.100000n V_hig
+ 432.100001n V_hig
+ 432.200000n V_hig
+ 432.200001n V_hig
+ 432.300000n V_hig
+ 432.300001n V_hig
+ 432.400000n V_hig
+ 432.400001n V_hig
+ 432.500000n V_hig
+ 432.500001n V_hig
+ 432.600000n V_hig
+ 432.600001n V_hig
+ 432.700000n V_hig
+ 432.700001n V_hig
+ 432.800000n V_hig
+ 432.800001n V_hig
+ 432.900000n V_hig
+ 432.900001n V_hig
+ 433.000000n V_hig
+ 433.000001n V_hig
+ 433.100000n V_hig
+ 433.100001n V_hig
+ 433.200000n V_hig
+ 433.200001n V_hig
+ 433.300000n V_hig
+ 433.300001n V_hig
+ 433.400000n V_hig
+ 433.400001n V_hig
+ 433.500000n V_hig
+ 433.500001n V_hig
+ 433.600000n V_hig
+ 433.600001n V_hig
+ 433.700000n V_hig
+ 433.700001n V_hig
+ 433.800000n V_hig
+ 433.800001n V_hig
+ 433.900000n V_hig
+ 433.900001n V_hig
+ 434.000000n V_hig
+ 434.000001n V_low
+ 434.100000n V_low
+ 434.100001n V_low
+ 434.200000n V_low
+ 434.200001n V_low
+ 434.300000n V_low
+ 434.300001n V_low
+ 434.400000n V_low
+ 434.400001n V_low
+ 434.500000n V_low
+ 434.500001n V_low
+ 434.600000n V_low
+ 434.600001n V_low
+ 434.700000n V_low
+ 434.700001n V_low
+ 434.800000n V_low
+ 434.800001n V_low
+ 434.900000n V_low
+ 434.900001n V_low
+ 435.000000n V_low
+ 435.000001n V_low
+ 435.100000n V_low
+ 435.100001n V_low
+ 435.200000n V_low
+ 435.200001n V_low
+ 435.300000n V_low
+ 435.300001n V_low
+ 435.400000n V_low
+ 435.400001n V_low
+ 435.500000n V_low
+ 435.500001n V_low
+ 435.600000n V_low
+ 435.600001n V_low
+ 435.700000n V_low
+ 435.700001n V_low
+ 435.800000n V_low
+ 435.800001n V_low
+ 435.900000n V_low
+ 435.900001n V_low
+ 436.000000n V_low
+ 436.000001n V_low
+ 436.100000n V_low
+ 436.100001n V_low
+ 436.200000n V_low
+ 436.200001n V_low
+ 436.300000n V_low
+ 436.300001n V_low
+ 436.400000n V_low
+ 436.400001n V_low
+ 436.500000n V_low
+ 436.500001n V_low
+ 436.600000n V_low
+ 436.600001n V_low
+ 436.700000n V_low
+ 436.700001n V_low
+ 436.800000n V_low
+ 436.800001n V_low
+ 436.900000n V_low
+ 436.900001n V_low
+ 437.000000n V_low
+ 437.000001n V_low
+ 437.100000n V_low
+ 437.100001n V_low
+ 437.200000n V_low
+ 437.200001n V_low
+ 437.300000n V_low
+ 437.300001n V_low
+ 437.400000n V_low
+ 437.400001n V_low
+ 437.500000n V_low
+ 437.500001n V_low
+ 437.600000n V_low
+ 437.600001n V_low
+ 437.700000n V_low
+ 437.700001n V_low
+ 437.800000n V_low
+ 437.800001n V_low
+ 437.900000n V_low
+ 437.900001n V_low
+ 438.000000n V_low
+ 438.000001n V_low
+ 438.100000n V_low
+ 438.100001n V_low
+ 438.200000n V_low
+ 438.200001n V_low
+ 438.300000n V_low
+ 438.300001n V_low
+ 438.400000n V_low
+ 438.400001n V_low
+ 438.500000n V_low
+ 438.500001n V_low
+ 438.600000n V_low
+ 438.600001n V_low
+ 438.700000n V_low
+ 438.700001n V_low
+ 438.800000n V_low
+ 438.800001n V_low
+ 438.900000n V_low
+ 438.900001n V_low
+ 439.000000n V_low
+ 439.000001n V_low
+ 439.100000n V_low
+ 439.100001n V_low
+ 439.200000n V_low
+ 439.200001n V_low
+ 439.300000n V_low
+ 439.300001n V_low
+ 439.400000n V_low
+ 439.400001n V_low
+ 439.500000n V_low
+ 439.500001n V_low
+ 439.600000n V_low
+ 439.600001n V_low
+ 439.700000n V_low
+ 439.700001n V_low
+ 439.800000n V_low
+ 439.800001n V_low
+ 439.900000n V_low
+ 439.900001n V_low
+ 440.000000n V_low
+ 440.000001n V_hig
+ 440.100000n V_hig
+ 440.100001n V_hig
+ 440.200000n V_hig
+ 440.200001n V_hig
+ 440.300000n V_hig
+ 440.300001n V_hig
+ 440.400000n V_hig
+ 440.400001n V_hig
+ 440.500000n V_hig
+ 440.500001n V_hig
+ 440.600000n V_hig
+ 440.600001n V_hig
+ 440.700000n V_hig
+ 440.700001n V_hig
+ 440.800000n V_hig
+ 440.800001n V_hig
+ 440.900000n V_hig
+ 440.900001n V_hig
+ 441.000000n V_hig
+ 441.000001n V_hig
+ 441.100000n V_hig
+ 441.100001n V_hig
+ 441.200000n V_hig
+ 441.200001n V_hig
+ 441.300000n V_hig
+ 441.300001n V_hig
+ 441.400000n V_hig
+ 441.400001n V_hig
+ 441.500000n V_hig
+ 441.500001n V_hig
+ 441.600000n V_hig
+ 441.600001n V_hig
+ 441.700000n V_hig
+ 441.700001n V_hig
+ 441.800000n V_hig
+ 441.800001n V_hig
+ 441.900000n V_hig
+ 441.900001n V_hig
+ 442.000000n V_hig
+ 442.000001n V_hig
+ 442.100000n V_hig
+ 442.100001n V_hig
+ 442.200000n V_hig
+ 442.200001n V_hig
+ 442.300000n V_hig
+ 442.300001n V_hig
+ 442.400000n V_hig
+ 442.400001n V_hig
+ 442.500000n V_hig
+ 442.500001n V_hig
+ 442.600000n V_hig
+ 442.600001n V_hig
+ 442.700000n V_hig
+ 442.700001n V_hig
+ 442.800000n V_hig
+ 442.800001n V_hig
+ 442.900000n V_hig
+ 442.900001n V_hig
+ 443.000000n V_hig
+ 443.000001n V_hig
+ 443.100000n V_hig
+ 443.100001n V_hig
+ 443.200000n V_hig
+ 443.200001n V_hig
+ 443.300000n V_hig
+ 443.300001n V_hig
+ 443.400000n V_hig
+ 443.400001n V_hig
+ 443.500000n V_hig
+ 443.500001n V_hig
+ 443.600000n V_hig
+ 443.600001n V_hig
+ 443.700000n V_hig
+ 443.700001n V_hig
+ 443.800000n V_hig
+ 443.800001n V_hig
+ 443.900000n V_hig
+ 443.900001n V_hig
+ 444.000000n V_hig
+ 444.000001n V_hig
+ 444.100000n V_hig
+ 444.100001n V_hig
+ 444.200000n V_hig
+ 444.200001n V_hig
+ 444.300000n V_hig
+ 444.300001n V_hig
+ 444.400000n V_hig
+ 444.400001n V_hig
+ 444.500000n V_hig
+ 444.500001n V_hig
+ 444.600000n V_hig
+ 444.600001n V_hig
+ 444.700000n V_hig
+ 444.700001n V_hig
+ 444.800000n V_hig
+ 444.800001n V_hig
+ 444.900000n V_hig
+ 444.900001n V_hig
+ 445.000000n V_hig
+ 445.000001n V_low
+ 445.100000n V_low
+ 445.100001n V_low
+ 445.200000n V_low
+ 445.200001n V_low
+ 445.300000n V_low
+ 445.300001n V_low
+ 445.400000n V_low
+ 445.400001n V_low
+ 445.500000n V_low
+ 445.500001n V_low
+ 445.600000n V_low
+ 445.600001n V_low
+ 445.700000n V_low
+ 445.700001n V_low
+ 445.800000n V_low
+ 445.800001n V_low
+ 445.900000n V_low
+ 445.900001n V_low
+ 446.000000n V_low
+ 446.000001n V_hig
+ 446.100000n V_hig
+ 446.100001n V_hig
+ 446.200000n V_hig
+ 446.200001n V_hig
+ 446.300000n V_hig
+ 446.300001n V_hig
+ 446.400000n V_hig
+ 446.400001n V_hig
+ 446.500000n V_hig
+ 446.500001n V_hig
+ 446.600000n V_hig
+ 446.600001n V_hig
+ 446.700000n V_hig
+ 446.700001n V_hig
+ 446.800000n V_hig
+ 446.800001n V_hig
+ 446.900000n V_hig
+ 446.900001n V_hig
+ 447.000000n V_hig
+ 447.000001n V_low
+ 447.100000n V_low
+ 447.100001n V_low
+ 447.200000n V_low
+ 447.200001n V_low
+ 447.300000n V_low
+ 447.300001n V_low
+ 447.400000n V_low
+ 447.400001n V_low
+ 447.500000n V_low
+ 447.500001n V_low
+ 447.600000n V_low
+ 447.600001n V_low
+ 447.700000n V_low
+ 447.700001n V_low
+ 447.800000n V_low
+ 447.800001n V_low
+ 447.900000n V_low
+ 447.900001n V_low
+ 448.000000n V_low
+ 448.000001n V_low
+ 448.100000n V_low
+ 448.100001n V_low
+ 448.200000n V_low
+ 448.200001n V_low
+ 448.300000n V_low
+ 448.300001n V_low
+ 448.400000n V_low
+ 448.400001n V_low
+ 448.500000n V_low
+ 448.500001n V_low
+ 448.600000n V_low
+ 448.600001n V_low
+ 448.700000n V_low
+ 448.700001n V_low
+ 448.800000n V_low
+ 448.800001n V_low
+ 448.900000n V_low
+ 448.900001n V_low
+ 449.000000n V_low
+ 449.000001n V_hig
+ 449.100000n V_hig
+ 449.100001n V_hig
+ 449.200000n V_hig
+ 449.200001n V_hig
+ 449.300000n V_hig
+ 449.300001n V_hig
+ 449.400000n V_hig
+ 449.400001n V_hig
+ 449.500000n V_hig
+ 449.500001n V_hig
+ 449.600000n V_hig
+ 449.600001n V_hig
+ 449.700000n V_hig
+ 449.700001n V_hig
+ 449.800000n V_hig
+ 449.800001n V_hig
+ 449.900000n V_hig
+ 449.900001n V_hig
+ 450.000000n V_hig
+ 450.000001n V_hig
+ 450.100000n V_hig
+ 450.100001n V_hig
+ 450.200000n V_hig
+ 450.200001n V_hig
+ 450.300000n V_hig
+ 450.300001n V_hig
+ 450.400000n V_hig
+ 450.400001n V_hig
+ 450.500000n V_hig
+ 450.500001n V_hig
+ 450.600000n V_hig
+ 450.600001n V_hig
+ 450.700000n V_hig
+ 450.700001n V_hig
+ 450.800000n V_hig
+ 450.800001n V_hig
+ 450.900000n V_hig
+ 450.900001n V_hig
+ 451.000000n V_hig
+ 451.000001n V_low
+ 451.100000n V_low
+ 451.100001n V_low
+ 451.200000n V_low
+ 451.200001n V_low
+ 451.300000n V_low
+ 451.300001n V_low
+ 451.400000n V_low
+ 451.400001n V_low
+ 451.500000n V_low
+ 451.500001n V_low
+ 451.600000n V_low
+ 451.600001n V_low
+ 451.700000n V_low
+ 451.700001n V_low
+ 451.800000n V_low
+ 451.800001n V_low
+ 451.900000n V_low
+ 451.900001n V_low
+ 452.000000n V_low
+ 452.000001n V_low
+ 452.100000n V_low
+ 452.100001n V_low
+ 452.200000n V_low
+ 452.200001n V_low
+ 452.300000n V_low
+ 452.300001n V_low
+ 452.400000n V_low
+ 452.400001n V_low
+ 452.500000n V_low
+ 452.500001n V_low
+ 452.600000n V_low
+ 452.600001n V_low
+ 452.700000n V_low
+ 452.700001n V_low
+ 452.800000n V_low
+ 452.800001n V_low
+ 452.900000n V_low
+ 452.900001n V_low
+ 453.000000n V_low
+ 453.000001n V_low
+ 453.100000n V_low
+ 453.100001n V_low
+ 453.200000n V_low
+ 453.200001n V_low
+ 453.300000n V_low
+ 453.300001n V_low
+ 453.400000n V_low
+ 453.400001n V_low
+ 453.500000n V_low
+ 453.500001n V_low
+ 453.600000n V_low
+ 453.600001n V_low
+ 453.700000n V_low
+ 453.700001n V_low
+ 453.800000n V_low
+ 453.800001n V_low
+ 453.900000n V_low
+ 453.900001n V_low
+ 454.000000n V_low
+ 454.000001n V_hig
+ 454.100000n V_hig
+ 454.100001n V_hig
+ 454.200000n V_hig
+ 454.200001n V_hig
+ 454.300000n V_hig
+ 454.300001n V_hig
+ 454.400000n V_hig
+ 454.400001n V_hig
+ 454.500000n V_hig
+ 454.500001n V_hig
+ 454.600000n V_hig
+ 454.600001n V_hig
+ 454.700000n V_hig
+ 454.700001n V_hig
+ 454.800000n V_hig
+ 454.800001n V_hig
+ 454.900000n V_hig
+ 454.900001n V_hig
+ 455.000000n V_hig
+ 455.000001n V_low
+ 455.100000n V_low
+ 455.100001n V_low
+ 455.200000n V_low
+ 455.200001n V_low
+ 455.300000n V_low
+ 455.300001n V_low
+ 455.400000n V_low
+ 455.400001n V_low
+ 455.500000n V_low
+ 455.500001n V_low
+ 455.600000n V_low
+ 455.600001n V_low
+ 455.700000n V_low
+ 455.700001n V_low
+ 455.800000n V_low
+ 455.800001n V_low
+ 455.900000n V_low
+ 455.900001n V_low
+ 456.000000n V_low
+ 456.000001n V_low
+ 456.100000n V_low
+ 456.100001n V_low
+ 456.200000n V_low
+ 456.200001n V_low
+ 456.300000n V_low
+ 456.300001n V_low
+ 456.400000n V_low
+ 456.400001n V_low
+ 456.500000n V_low
+ 456.500001n V_low
+ 456.600000n V_low
+ 456.600001n V_low
+ 456.700000n V_low
+ 456.700001n V_low
+ 456.800000n V_low
+ 456.800001n V_low
+ 456.900000n V_low
+ 456.900001n V_low
+ 457.000000n V_low
+ 457.000001n V_hig
+ 457.100000n V_hig
+ 457.100001n V_hig
+ 457.200000n V_hig
+ 457.200001n V_hig
+ 457.300000n V_hig
+ 457.300001n V_hig
+ 457.400000n V_hig
+ 457.400001n V_hig
+ 457.500000n V_hig
+ 457.500001n V_hig
+ 457.600000n V_hig
+ 457.600001n V_hig
+ 457.700000n V_hig
+ 457.700001n V_hig
+ 457.800000n V_hig
+ 457.800001n V_hig
+ 457.900000n V_hig
+ 457.900001n V_hig
+ 458.000000n V_hig
+ 458.000001n V_hig
+ 458.100000n V_hig
+ 458.100001n V_hig
+ 458.200000n V_hig
+ 458.200001n V_hig
+ 458.300000n V_hig
+ 458.300001n V_hig
+ 458.400000n V_hig
+ 458.400001n V_hig
+ 458.500000n V_hig
+ 458.500001n V_hig
+ 458.600000n V_hig
+ 458.600001n V_hig
+ 458.700000n V_hig
+ 458.700001n V_hig
+ 458.800000n V_hig
+ 458.800001n V_hig
+ 458.900000n V_hig
+ 458.900001n V_hig
+ 459.000000n V_hig
+ 459.000001n V_low
+ 459.100000n V_low
+ 459.100001n V_low
+ 459.200000n V_low
+ 459.200001n V_low
+ 459.300000n V_low
+ 459.300001n V_low
+ 459.400000n V_low
+ 459.400001n V_low
+ 459.500000n V_low
+ 459.500001n V_low
+ 459.600000n V_low
+ 459.600001n V_low
+ 459.700000n V_low
+ 459.700001n V_low
+ 459.800000n V_low
+ 459.800001n V_low
+ 459.900000n V_low
+ 459.900001n V_low
+ 460.000000n V_low
+ 460.000001n V_hig
+ 460.100000n V_hig
+ 460.100001n V_hig
+ 460.200000n V_hig
+ 460.200001n V_hig
+ 460.300000n V_hig
+ 460.300001n V_hig
+ 460.400000n V_hig
+ 460.400001n V_hig
+ 460.500000n V_hig
+ 460.500001n V_hig
+ 460.600000n V_hig
+ 460.600001n V_hig
+ 460.700000n V_hig
+ 460.700001n V_hig
+ 460.800000n V_hig
+ 460.800001n V_hig
+ 460.900000n V_hig
+ 460.900001n V_hig
+ 461.000000n V_hig
+ 461.000001n V_low
+ 461.100000n V_low
+ 461.100001n V_low
+ 461.200000n V_low
+ 461.200001n V_low
+ 461.300000n V_low
+ 461.300001n V_low
+ 461.400000n V_low
+ 461.400001n V_low
+ 461.500000n V_low
+ 461.500001n V_low
+ 461.600000n V_low
+ 461.600001n V_low
+ 461.700000n V_low
+ 461.700001n V_low
+ 461.800000n V_low
+ 461.800001n V_low
+ 461.900000n V_low
+ 461.900001n V_low
+ 462.000000n V_low
+ 462.000001n V_low
+ 462.100000n V_low
+ 462.100001n V_low
+ 462.200000n V_low
+ 462.200001n V_low
+ 462.300000n V_low
+ 462.300001n V_low
+ 462.400000n V_low
+ 462.400001n V_low
+ 462.500000n V_low
+ 462.500001n V_low
+ 462.600000n V_low
+ 462.600001n V_low
+ 462.700000n V_low
+ 462.700001n V_low
+ 462.800000n V_low
+ 462.800001n V_low
+ 462.900000n V_low
+ 462.900001n V_low
+ 463.000000n V_low
+ 463.000001n V_low
+ 463.100000n V_low
+ 463.100001n V_low
+ 463.200000n V_low
+ 463.200001n V_low
+ 463.300000n V_low
+ 463.300001n V_low
+ 463.400000n V_low
+ 463.400001n V_low
+ 463.500000n V_low
+ 463.500001n V_low
+ 463.600000n V_low
+ 463.600001n V_low
+ 463.700000n V_low
+ 463.700001n V_low
+ 463.800000n V_low
+ 463.800001n V_low
+ 463.900000n V_low
+ 463.900001n V_low
+ 464.000000n V_low
+ 464.000001n V_hig
+ 464.100000n V_hig
+ 464.100001n V_hig
+ 464.200000n V_hig
+ 464.200001n V_hig
+ 464.300000n V_hig
+ 464.300001n V_hig
+ 464.400000n V_hig
+ 464.400001n V_hig
+ 464.500000n V_hig
+ 464.500001n V_hig
+ 464.600000n V_hig
+ 464.600001n V_hig
+ 464.700000n V_hig
+ 464.700001n V_hig
+ 464.800000n V_hig
+ 464.800001n V_hig
+ 464.900000n V_hig
+ 464.900001n V_hig
+ 465.000000n V_hig
+ 465.000001n V_low
+ 465.100000n V_low
+ 465.100001n V_low
+ 465.200000n V_low
+ 465.200001n V_low
+ 465.300000n V_low
+ 465.300001n V_low
+ 465.400000n V_low
+ 465.400001n V_low
+ 465.500000n V_low
+ 465.500001n V_low
+ 465.600000n V_low
+ 465.600001n V_low
+ 465.700000n V_low
+ 465.700001n V_low
+ 465.800000n V_low
+ 465.800001n V_low
+ 465.900000n V_low
+ 465.900001n V_low
+ 466.000000n V_low
+ 466.000001n V_low
+ 466.100000n V_low
+ 466.100001n V_low
+ 466.200000n V_low
+ 466.200001n V_low
+ 466.300000n V_low
+ 466.300001n V_low
+ 466.400000n V_low
+ 466.400001n V_low
+ 466.500000n V_low
+ 466.500001n V_low
+ 466.600000n V_low
+ 466.600001n V_low
+ 466.700000n V_low
+ 466.700001n V_low
+ 466.800000n V_low
+ 466.800001n V_low
+ 466.900000n V_low
+ 466.900001n V_low
+ 467.000000n V_low
+ 467.000001n V_low
+ 467.100000n V_low
+ 467.100001n V_low
+ 467.200000n V_low
+ 467.200001n V_low
+ 467.300000n V_low
+ 467.300001n V_low
+ 467.400000n V_low
+ 467.400001n V_low
+ 467.500000n V_low
+ 467.500001n V_low
+ 467.600000n V_low
+ 467.600001n V_low
+ 467.700000n V_low
+ 467.700001n V_low
+ 467.800000n V_low
+ 467.800001n V_low
+ 467.900000n V_low
+ 467.900001n V_low
+ 468.000000n V_low
+ 468.000001n V_hig
+ 468.100000n V_hig
+ 468.100001n V_hig
+ 468.200000n V_hig
+ 468.200001n V_hig
+ 468.300000n V_hig
+ 468.300001n V_hig
+ 468.400000n V_hig
+ 468.400001n V_hig
+ 468.500000n V_hig
+ 468.500001n V_hig
+ 468.600000n V_hig
+ 468.600001n V_hig
+ 468.700000n V_hig
+ 468.700001n V_hig
+ 468.800000n V_hig
+ 468.800001n V_hig
+ 468.900000n V_hig
+ 468.900001n V_hig
+ 469.000000n V_hig
+ 469.000001n V_low
+ 469.100000n V_low
+ 469.100001n V_low
+ 469.200000n V_low
+ 469.200001n V_low
+ 469.300000n V_low
+ 469.300001n V_low
+ 469.400000n V_low
+ 469.400001n V_low
+ 469.500000n V_low
+ 469.500001n V_low
+ 469.600000n V_low
+ 469.600001n V_low
+ 469.700000n V_low
+ 469.700001n V_low
+ 469.800000n V_low
+ 469.800001n V_low
+ 469.900000n V_low
+ 469.900001n V_low
+ 470.000000n V_low
+ 470.000001n V_low
+ 470.100000n V_low
+ 470.100001n V_low
+ 470.200000n V_low
+ 470.200001n V_low
+ 470.300000n V_low
+ 470.300001n V_low
+ 470.400000n V_low
+ 470.400001n V_low
+ 470.500000n V_low
+ 470.500001n V_low
+ 470.600000n V_low
+ 470.600001n V_low
+ 470.700000n V_low
+ 470.700001n V_low
+ 470.800000n V_low
+ 470.800001n V_low
+ 470.900000n V_low
+ 470.900001n V_low
+ 471.000000n V_low
+ 471.000001n V_hig
+ 471.100000n V_hig
+ 471.100001n V_hig
+ 471.200000n V_hig
+ 471.200001n V_hig
+ 471.300000n V_hig
+ 471.300001n V_hig
+ 471.400000n V_hig
+ 471.400001n V_hig
+ 471.500000n V_hig
+ 471.500001n V_hig
+ 471.600000n V_hig
+ 471.600001n V_hig
+ 471.700000n V_hig
+ 471.700001n V_hig
+ 471.800000n V_hig
+ 471.800001n V_hig
+ 471.900000n V_hig
+ 471.900001n V_hig
+ 472.000000n V_hig
+ 472.000001n V_low
+ 472.100000n V_low
+ 472.100001n V_low
+ 472.200000n V_low
+ 472.200001n V_low
+ 472.300000n V_low
+ 472.300001n V_low
+ 472.400000n V_low
+ 472.400001n V_low
+ 472.500000n V_low
+ 472.500001n V_low
+ 472.600000n V_low
+ 472.600001n V_low
+ 472.700000n V_low
+ 472.700001n V_low
+ 472.800000n V_low
+ 472.800001n V_low
+ 472.900000n V_low
+ 472.900001n V_low
+ 473.000000n V_low
+ 473.000001n V_low
+ 473.100000n V_low
+ 473.100001n V_low
+ 473.200000n V_low
+ 473.200001n V_low
+ 473.300000n V_low
+ 473.300001n V_low
+ 473.400000n V_low
+ 473.400001n V_low
+ 473.500000n V_low
+ 473.500001n V_low
+ 473.600000n V_low
+ 473.600001n V_low
+ 473.700000n V_low
+ 473.700001n V_low
+ 473.800000n V_low
+ 473.800001n V_low
+ 473.900000n V_low
+ 473.900001n V_low
+ 474.000000n V_low
+ 474.000001n V_low
+ 474.100000n V_low
+ 474.100001n V_low
+ 474.200000n V_low
+ 474.200001n V_low
+ 474.300000n V_low
+ 474.300001n V_low
+ 474.400000n V_low
+ 474.400001n V_low
+ 474.500000n V_low
+ 474.500001n V_low
+ 474.600000n V_low
+ 474.600001n V_low
+ 474.700000n V_low
+ 474.700001n V_low
+ 474.800000n V_low
+ 474.800001n V_low
+ 474.900000n V_low
+ 474.900001n V_low
+ 475.000000n V_low
+ 475.000001n V_hig
+ 475.100000n V_hig
+ 475.100001n V_hig
+ 475.200000n V_hig
+ 475.200001n V_hig
+ 475.300000n V_hig
+ 475.300001n V_hig
+ 475.400000n V_hig
+ 475.400001n V_hig
+ 475.500000n V_hig
+ 475.500001n V_hig
+ 475.600000n V_hig
+ 475.600001n V_hig
+ 475.700000n V_hig
+ 475.700001n V_hig
+ 475.800000n V_hig
+ 475.800001n V_hig
+ 475.900000n V_hig
+ 475.900001n V_hig
+ 476.000000n V_hig
+ 476.000001n V_hig
+ 476.100000n V_hig
+ 476.100001n V_hig
+ 476.200000n V_hig
+ 476.200001n V_hig
+ 476.300000n V_hig
+ 476.300001n V_hig
+ 476.400000n V_hig
+ 476.400001n V_hig
+ 476.500000n V_hig
+ 476.500001n V_hig
+ 476.600000n V_hig
+ 476.600001n V_hig
+ 476.700000n V_hig
+ 476.700001n V_hig
+ 476.800000n V_hig
+ 476.800001n V_hig
+ 476.900000n V_hig
+ 476.900001n V_hig
+ 477.000000n V_hig
+ 477.000001n V_low
+ 477.100000n V_low
+ 477.100001n V_low
+ 477.200000n V_low
+ 477.200001n V_low
+ 477.300000n V_low
+ 477.300001n V_low
+ 477.400000n V_low
+ 477.400001n V_low
+ 477.500000n V_low
+ 477.500001n V_low
+ 477.600000n V_low
+ 477.600001n V_low
+ 477.700000n V_low
+ 477.700001n V_low
+ 477.800000n V_low
+ 477.800001n V_low
+ 477.900000n V_low
+ 477.900001n V_low
+ 478.000000n V_low
+ 478.000001n V_hig
+ 478.100000n V_hig
+ 478.100001n V_hig
+ 478.200000n V_hig
+ 478.200001n V_hig
+ 478.300000n V_hig
+ 478.300001n V_hig
+ 478.400000n V_hig
+ 478.400001n V_hig
+ 478.500000n V_hig
+ 478.500001n V_hig
+ 478.600000n V_hig
+ 478.600001n V_hig
+ 478.700000n V_hig
+ 478.700001n V_hig
+ 478.800000n V_hig
+ 478.800001n V_hig
+ 478.900000n V_hig
+ 478.900001n V_hig
+ 479.000000n V_hig
+ 479.000001n V_hig
+ 479.100000n V_hig
+ 479.100001n V_hig
+ 479.200000n V_hig
+ 479.200001n V_hig
+ 479.300000n V_hig
+ 479.300001n V_hig
+ 479.400000n V_hig
+ 479.400001n V_hig
+ 479.500000n V_hig
+ 479.500001n V_hig
+ 479.600000n V_hig
+ 479.600001n V_hig
+ 479.700000n V_hig
+ 479.700001n V_hig
+ 479.800000n V_hig
+ 479.800001n V_hig
+ 479.900000n V_hig
+ 479.900001n V_hig
+ 480.000000n V_hig
+ 480.000001n V_hig
+ 480.100000n V_hig
+ 480.100001n V_hig
+ 480.200000n V_hig
+ 480.200001n V_hig
+ 480.300000n V_hig
+ 480.300001n V_hig
+ 480.400000n V_hig
+ 480.400001n V_hig
+ 480.500000n V_hig
+ 480.500001n V_hig
+ 480.600000n V_hig
+ 480.600001n V_hig
+ 480.700000n V_hig
+ 480.700001n V_hig
+ 480.800000n V_hig
+ 480.800001n V_hig
+ 480.900000n V_hig
+ 480.900001n V_hig
+ 481.000000n V_hig
+ 481.000001n V_hig
+ 481.100000n V_hig
+ 481.100001n V_hig
+ 481.200000n V_hig
+ 481.200001n V_hig
+ 481.300000n V_hig
+ 481.300001n V_hig
+ 481.400000n V_hig
+ 481.400001n V_hig
+ 481.500000n V_hig
+ 481.500001n V_hig
+ 481.600000n V_hig
+ 481.600001n V_hig
+ 481.700000n V_hig
+ 481.700001n V_hig
+ 481.800000n V_hig
+ 481.800001n V_hig
+ 481.900000n V_hig
+ 481.900001n V_hig
+ 482.000000n V_hig
+ 482.000001n V_low
+ 482.100000n V_low
+ 482.100001n V_low
+ 482.200000n V_low
+ 482.200001n V_low
+ 482.300000n V_low
+ 482.300001n V_low
+ 482.400000n V_low
+ 482.400001n V_low
+ 482.500000n V_low
+ 482.500001n V_low
+ 482.600000n V_low
+ 482.600001n V_low
+ 482.700000n V_low
+ 482.700001n V_low
+ 482.800000n V_low
+ 482.800001n V_low
+ 482.900000n V_low
+ 482.900001n V_low
+ 483.000000n V_low
+ 483.000001n V_low
+ 483.100000n V_low
+ 483.100001n V_low
+ 483.200000n V_low
+ 483.200001n V_low
+ 483.300000n V_low
+ 483.300001n V_low
+ 483.400000n V_low
+ 483.400001n V_low
+ 483.500000n V_low
+ 483.500001n V_low
+ 483.600000n V_low
+ 483.600001n V_low
+ 483.700000n V_low
+ 483.700001n V_low
+ 483.800000n V_low
+ 483.800001n V_low
+ 483.900000n V_low
+ 483.900001n V_low
+ 484.000000n V_low
+ 484.000001n V_low
+ 484.100000n V_low
+ 484.100001n V_low
+ 484.200000n V_low
+ 484.200001n V_low
+ 484.300000n V_low
+ 484.300001n V_low
+ 484.400000n V_low
+ 484.400001n V_low
+ 484.500000n V_low
+ 484.500001n V_low
+ 484.600000n V_low
+ 484.600001n V_low
+ 484.700000n V_low
+ 484.700001n V_low
+ 484.800000n V_low
+ 484.800001n V_low
+ 484.900000n V_low
+ 484.900001n V_low
+ 485.000000n V_low
+ 485.000001n V_low
+ 485.100000n V_low
+ 485.100001n V_low
+ 485.200000n V_low
+ 485.200001n V_low
+ 485.300000n V_low
+ 485.300001n V_low
+ 485.400000n V_low
+ 485.400001n V_low
+ 485.500000n V_low
+ 485.500001n V_low
+ 485.600000n V_low
+ 485.600001n V_low
+ 485.700000n V_low
+ 485.700001n V_low
+ 485.800000n V_low
+ 485.800001n V_low
+ 485.900000n V_low
+ 485.900001n V_low
+ 486.000000n V_low
+ 486.000001n V_low
+ 486.100000n V_low
+ 486.100001n V_low
+ 486.200000n V_low
+ 486.200001n V_low
+ 486.300000n V_low
+ 486.300001n V_low
+ 486.400000n V_low
+ 486.400001n V_low
+ 486.500000n V_low
+ 486.500001n V_low
+ 486.600000n V_low
+ 486.600001n V_low
+ 486.700000n V_low
+ 486.700001n V_low
+ 486.800000n V_low
+ 486.800001n V_low
+ 486.900000n V_low
+ 486.900001n V_low
+ 487.000000n V_low
+ 487.000001n V_low
+ 487.100000n V_low
+ 487.100001n V_low
+ 487.200000n V_low
+ 487.200001n V_low
+ 487.300000n V_low
+ 487.300001n V_low
+ 487.400000n V_low
+ 487.400001n V_low
+ 487.500000n V_low
+ 487.500001n V_low
+ 487.600000n V_low
+ 487.600001n V_low
+ 487.700000n V_low
+ 487.700001n V_low
+ 487.800000n V_low
+ 487.800001n V_low
+ 487.900000n V_low
+ 487.900001n V_low
+ 488.000000n V_low
+ 488.000001n V_hig
+ 488.100000n V_hig
+ 488.100001n V_hig
+ 488.200000n V_hig
+ 488.200001n V_hig
+ 488.300000n V_hig
+ 488.300001n V_hig
+ 488.400000n V_hig
+ 488.400001n V_hig
+ 488.500000n V_hig
+ 488.500001n V_hig
+ 488.600000n V_hig
+ 488.600001n V_hig
+ 488.700000n V_hig
+ 488.700001n V_hig
+ 488.800000n V_hig
+ 488.800001n V_hig
+ 488.900000n V_hig
+ 488.900001n V_hig
+ 489.000000n V_hig
+ 489.000001n V_hig
+ 489.100000n V_hig
+ 489.100001n V_hig
+ 489.200000n V_hig
+ 489.200001n V_hig
+ 489.300000n V_hig
+ 489.300001n V_hig
+ 489.400000n V_hig
+ 489.400001n V_hig
+ 489.500000n V_hig
+ 489.500001n V_hig
+ 489.600000n V_hig
+ 489.600001n V_hig
+ 489.700000n V_hig
+ 489.700001n V_hig
+ 489.800000n V_hig
+ 489.800001n V_hig
+ 489.900000n V_hig
+ 489.900001n V_hig
+ 490.000000n V_hig
+ 490.000001n V_hig
+ 490.100000n V_hig
+ 490.100001n V_hig
+ 490.200000n V_hig
+ 490.200001n V_hig
+ 490.300000n V_hig
+ 490.300001n V_hig
+ 490.400000n V_hig
+ 490.400001n V_hig
+ 490.500000n V_hig
+ 490.500001n V_hig
+ 490.600000n V_hig
+ 490.600001n V_hig
+ 490.700000n V_hig
+ 490.700001n V_hig
+ 490.800000n V_hig
+ 490.800001n V_hig
+ 490.900000n V_hig
+ 490.900001n V_hig
+ 491.000000n V_hig
+ 491.000001n V_hig
+ 491.100000n V_hig
+ 491.100001n V_hig
+ 491.200000n V_hig
+ 491.200001n V_hig
+ 491.300000n V_hig
+ 491.300001n V_hig
+ 491.400000n V_hig
+ 491.400001n V_hig
+ 491.500000n V_hig
+ 491.500001n V_hig
+ 491.600000n V_hig
+ 491.600001n V_hig
+ 491.700000n V_hig
+ 491.700001n V_hig
+ 491.800000n V_hig
+ 491.800001n V_hig
+ 491.900000n V_hig
+ 491.900001n V_hig
+ 492.000000n V_hig
+ 492.000001n V_low
+ 492.100000n V_low
+ 492.100001n V_low
+ 492.200000n V_low
+ 492.200001n V_low
+ 492.300000n V_low
+ 492.300001n V_low
+ 492.400000n V_low
+ 492.400001n V_low
+ 492.500000n V_low
+ 492.500001n V_low
+ 492.600000n V_low
+ 492.600001n V_low
+ 492.700000n V_low
+ 492.700001n V_low
+ 492.800000n V_low
+ 492.800001n V_low
+ 492.900000n V_low
+ 492.900001n V_low
+ 493.000000n V_low
+ 493.000001n V_low
+ 493.100000n V_low
+ 493.100001n V_low
+ 493.200000n V_low
+ 493.200001n V_low
+ 493.300000n V_low
+ 493.300001n V_low
+ 493.400000n V_low
+ 493.400001n V_low
+ 493.500000n V_low
+ 493.500001n V_low
+ 493.600000n V_low
+ 493.600001n V_low
+ 493.700000n V_low
+ 493.700001n V_low
+ 493.800000n V_low
+ 493.800001n V_low
+ 493.900000n V_low
+ 493.900001n V_low
+ 494.000000n V_low
+ 494.000001n V_low
+ 494.100000n V_low
+ 494.100001n V_low
+ 494.200000n V_low
+ 494.200001n V_low
+ 494.300000n V_low
+ 494.300001n V_low
+ 494.400000n V_low
+ 494.400001n V_low
+ 494.500000n V_low
+ 494.500001n V_low
+ 494.600000n V_low
+ 494.600001n V_low
+ 494.700000n V_low
+ 494.700001n V_low
+ 494.800000n V_low
+ 494.800001n V_low
+ 494.900000n V_low
+ 494.900001n V_low
+ 495.000000n V_low
+ 495.000001n V_hig
+ 495.100000n V_hig
+ 495.100001n V_hig
+ 495.200000n V_hig
+ 495.200001n V_hig
+ 495.300000n V_hig
+ 495.300001n V_hig
+ 495.400000n V_hig
+ 495.400001n V_hig
+ 495.500000n V_hig
+ 495.500001n V_hig
+ 495.600000n V_hig
+ 495.600001n V_hig
+ 495.700000n V_hig
+ 495.700001n V_hig
+ 495.800000n V_hig
+ 495.800001n V_hig
+ 495.900000n V_hig
+ 495.900001n V_hig
+ 496.000000n V_hig
+ 496.000001n V_hig
+ 496.100000n V_hig
+ 496.100001n V_hig
+ 496.200000n V_hig
+ 496.200001n V_hig
+ 496.300000n V_hig
+ 496.300001n V_hig
+ 496.400000n V_hig
+ 496.400001n V_hig
+ 496.500000n V_hig
+ 496.500001n V_hig
+ 496.600000n V_hig
+ 496.600001n V_hig
+ 496.700000n V_hig
+ 496.700001n V_hig
+ 496.800000n V_hig
+ 496.800001n V_hig
+ 496.900000n V_hig
+ 496.900001n V_hig
+ 497.000000n V_hig
+ 497.000001n V_hig
+ 497.100000n V_hig
+ 497.100001n V_hig
+ 497.200000n V_hig
+ 497.200001n V_hig
+ 497.300000n V_hig
+ 497.300001n V_hig
+ 497.400000n V_hig
+ 497.400001n V_hig
+ 497.500000n V_hig
+ 497.500001n V_hig
+ 497.600000n V_hig
+ 497.600001n V_hig
+ 497.700000n V_hig
+ 497.700001n V_hig
+ 497.800000n V_hig
+ 497.800001n V_hig
+ 497.900000n V_hig
+ 497.900001n V_hig
+ 498.000000n V_hig
+ 498.000001n V_hig
+ 498.100000n V_hig
+ 498.100001n V_hig
+ 498.200000n V_hig
+ 498.200001n V_hig
+ 498.300000n V_hig
+ 498.300001n V_hig
+ 498.400000n V_hig
+ 498.400001n V_hig
+ 498.500000n V_hig
+ 498.500001n V_hig
+ 498.600000n V_hig
+ 498.600001n V_hig
+ 498.700000n V_hig
+ 498.700001n V_hig
+ 498.800000n V_hig
+ 498.800001n V_hig
+ 498.900000n V_hig
+ 498.900001n V_hig
+ 499.000000n V_hig
+ 499.000001n V_hig
+ 499.100000n V_hig
+ 499.100001n V_hig
+ 499.200000n V_hig
+ 499.200001n V_hig
+ 499.300000n V_hig
+ 499.300001n V_hig
+ 499.400000n V_hig
+ 499.400001n V_hig
+ 499.500000n V_hig
+ 499.500001n V_hig
+ 499.600000n V_hig
+ 499.600001n V_hig
+ 499.700000n V_hig
+ 499.700001n V_hig
+ 499.800000n V_hig
+ 499.800001n V_hig
+ 499.900000n V_hig
+ 499.900001n V_hig
+ 500.000000n V_hig
+ 500.000001n V_low
+ 500.100000n V_low
+ 500.100001n V_low
+ 500.200000n V_low
+ 500.200001n V_low
+ 500.300000n V_low
+ 500.300001n V_low
+ 500.400000n V_low
+ 500.400001n V_low
+ 500.500000n V_low
+ 500.500001n V_low
+ 500.600000n V_low
+ 500.600001n V_low
+ 500.700000n V_low
+ 500.700001n V_low
+ 500.800000n V_low
+ 500.800001n V_low
+ 500.900000n V_low
+ 500.900001n V_low
+ 501.000000n V_low
+ 501.000001n V_low
+ 501.100000n V_low
+ 501.100001n V_low
+ 501.200000n V_low
+ 501.200001n V_low
+ 501.300000n V_low
+ 501.300001n V_low
+ 501.400000n V_low
+ 501.400001n V_low
+ 501.500000n V_low
+ 501.500001n V_low
+ 501.600000n V_low
+ 501.600001n V_low
+ 501.700000n V_low
+ 501.700001n V_low
+ 501.800000n V_low
+ 501.800001n V_low
+ 501.900000n V_low
+ 501.900001n V_low
+ 502.000000n V_low
+ 502.000001n V_low
+ 502.100000n V_low
+ 502.100001n V_low
+ 502.200000n V_low
+ 502.200001n V_low
+ 502.300000n V_low
+ 502.300001n V_low
+ 502.400000n V_low
+ 502.400001n V_low
+ 502.500000n V_low
+ 502.500001n V_low
+ 502.600000n V_low
+ 502.600001n V_low
+ 502.700000n V_low
+ 502.700001n V_low
+ 502.800000n V_low
+ 502.800001n V_low
+ 502.900000n V_low
+ 502.900001n V_low
+ 503.000000n V_low
+ 503.000001n V_low
+ 503.100000n V_low
+ 503.100001n V_low
+ 503.200000n V_low
+ 503.200001n V_low
+ 503.300000n V_low
+ 503.300001n V_low
+ 503.400000n V_low
+ 503.400001n V_low
+ 503.500000n V_low
+ 503.500001n V_low
+ 503.600000n V_low
+ 503.600001n V_low
+ 503.700000n V_low
+ 503.700001n V_low
+ 503.800000n V_low
+ 503.800001n V_low
+ 503.900000n V_low
+ 503.900001n V_low
+ 504.000000n V_low
+ 504.000001n V_low
+ 504.100000n V_low
+ 504.100001n V_low
+ 504.200000n V_low
+ 504.200001n V_low
+ 504.300000n V_low
+ 504.300001n V_low
+ 504.400000n V_low
+ 504.400001n V_low
+ 504.500000n V_low
+ 504.500001n V_low
+ 504.600000n V_low
+ 504.600001n V_low
+ 504.700000n V_low
+ 504.700001n V_low
+ 504.800000n V_low
+ 504.800001n V_low
+ 504.900000n V_low
+ 504.900001n V_low
+ 505.000000n V_low
+ 505.000001n V_low
+ 505.100000n V_low
+ 505.100001n V_low
+ 505.200000n V_low
+ 505.200001n V_low
+ 505.300000n V_low
+ 505.300001n V_low
+ 505.400000n V_low
+ 505.400001n V_low
+ 505.500000n V_low
+ 505.500001n V_low
+ 505.600000n V_low
+ 505.600001n V_low
+ 505.700000n V_low
+ 505.700001n V_low
+ 505.800000n V_low
+ 505.800001n V_low
+ 505.900000n V_low
+ 505.900001n V_low
+ 506.000000n V_low
+ 506.000001n V_low
+ 506.100000n V_low
+ 506.100001n V_low
+ 506.200000n V_low
+ 506.200001n V_low
+ 506.300000n V_low
+ 506.300001n V_low
+ 506.400000n V_low
+ 506.400001n V_low
+ 506.500000n V_low
+ 506.500001n V_low
+ 506.600000n V_low
+ 506.600001n V_low
+ 506.700000n V_low
+ 506.700001n V_low
+ 506.800000n V_low
+ 506.800001n V_low
+ 506.900000n V_low
+ 506.900001n V_low
+ 507.000000n V_low
+ 507.000001n V_hig
+ 507.100000n V_hig
+ 507.100001n V_hig
+ 507.200000n V_hig
+ 507.200001n V_hig
+ 507.300000n V_hig
+ 507.300001n V_hig
+ 507.400000n V_hig
+ 507.400001n V_hig
+ 507.500000n V_hig
+ 507.500001n V_hig
+ 507.600000n V_hig
+ 507.600001n V_hig
+ 507.700000n V_hig
+ 507.700001n V_hig
+ 507.800000n V_hig
+ 507.800001n V_hig
+ 507.900000n V_hig
+ 507.900001n V_hig
+ 508.000000n V_hig
+ 508.000001n V_low
+ 508.100000n V_low
+ 508.100001n V_low
+ 508.200000n V_low
+ 508.200001n V_low
+ 508.300000n V_low
+ 508.300001n V_low
+ 508.400000n V_low
+ 508.400001n V_low
+ 508.500000n V_low
+ 508.500001n V_low
+ 508.600000n V_low
+ 508.600001n V_low
+ 508.700000n V_low
+ 508.700001n V_low
+ 508.800000n V_low
+ 508.800001n V_low
+ 508.900000n V_low
+ 508.900001n V_low
+ 509.000000n V_low
+ 509.000001n V_hig
+ 509.100000n V_hig
+ 509.100001n V_hig
+ 509.200000n V_hig
+ 509.200001n V_hig
+ 509.300000n V_hig
+ 509.300001n V_hig
+ 509.400000n V_hig
+ 509.400001n V_hig
+ 509.500000n V_hig
+ 509.500001n V_hig
+ 509.600000n V_hig
+ 509.600001n V_hig
+ 509.700000n V_hig
+ 509.700001n V_hig
+ 509.800000n V_hig
+ 509.800001n V_hig
+ 509.900000n V_hig
+ 509.900001n V_hig
+ 510.000000n V_hig
+ 510.000001n V_hig
+ 510.100000n V_hig
+ 510.100001n V_hig
+ 510.200000n V_hig
+ 510.200001n V_hig
+ 510.300000n V_hig
+ 510.300001n V_hig
+ 510.400000n V_hig
+ 510.400001n V_hig
+ 510.500000n V_hig
+ 510.500001n V_hig
+ 510.600000n V_hig
+ 510.600001n V_hig
+ 510.700000n V_hig
+ 510.700001n V_hig
+ 510.800000n V_hig
+ 510.800001n V_hig
+ 510.900000n V_hig
+ 510.900001n V_hig
+ 511.000000n V_hig
+ 511.000001n V_hig
+ 511.100000n V_hig
+ 511.100001n V_hig
+ 511.200000n V_hig
+ 511.200001n V_hig
+ 511.300000n V_hig
+ 511.300001n V_hig
+ 511.400000n V_hig
+ 511.400001n V_hig
+ 511.500000n V_hig
+ 511.500001n V_hig
+ 511.600000n V_hig
+ 511.600001n V_hig
+ 511.700000n V_hig
+ 511.700001n V_hig
+ 511.800000n V_hig
+ 511.800001n V_hig
+ 511.900000n V_hig
+ 511.900001n V_hig
+ 512.000000n V_hig
+ 512.000001n V_hig
+ 512.100000n V_hig
+ 512.100001n V_hig
+ 512.200000n V_hig
+ 512.200001n V_hig
+ 512.300000n V_hig
+ 512.300001n V_hig
+ 512.400000n V_hig
+ 512.400001n V_hig
+ 512.500000n V_hig
+ 512.500001n V_hig
+ 512.600000n V_hig
+ 512.600001n V_hig
+ 512.700000n V_hig
+ 512.700001n V_hig
+ 512.800000n V_hig
+ 512.800001n V_hig
+ 512.900000n V_hig
+ 512.900001n V_hig
+ 513.000000n V_hig
+ 513.000001n V_low
+ 513.100000n V_low
+ 513.100001n V_low
+ 513.200000n V_low
+ 513.200001n V_low
+ 513.300000n V_low
+ 513.300001n V_low
+ 513.400000n V_low
+ 513.400001n V_low
+ 513.500000n V_low
+ 513.500001n V_low
+ 513.600000n V_low
+ 513.600001n V_low
+ 513.700000n V_low
+ 513.700001n V_low
+ 513.800000n V_low
+ 513.800001n V_low
+ 513.900000n V_low
+ 513.900001n V_low
+ 514.000000n V_low
+ 514.000001n V_low
+ 514.100000n V_low
+ 514.100001n V_low
+ 514.200000n V_low
+ 514.200001n V_low
+ 514.300000n V_low
+ 514.300001n V_low
+ 514.400000n V_low
+ 514.400001n V_low
+ 514.500000n V_low
+ 514.500001n V_low
+ 514.600000n V_low
+ 514.600001n V_low
+ 514.700000n V_low
+ 514.700001n V_low
+ 514.800000n V_low
+ 514.800001n V_low
+ 514.900000n V_low
+ 514.900001n V_low
+ 515.000000n V_low
+ 515.000001n V_hig
+ 515.100000n V_hig
+ 515.100001n V_hig
+ 515.200000n V_hig
+ 515.200001n V_hig
+ 515.300000n V_hig
+ 515.300001n V_hig
+ 515.400000n V_hig
+ 515.400001n V_hig
+ 515.500000n V_hig
+ 515.500001n V_hig
+ 515.600000n V_hig
+ 515.600001n V_hig
+ 515.700000n V_hig
+ 515.700001n V_hig
+ 515.800000n V_hig
+ 515.800001n V_hig
+ 515.900000n V_hig
+ 515.900001n V_hig
+ 516.000000n V_hig
+ 516.000001n V_low
+ 516.100000n V_low
+ 516.100001n V_low
+ 516.200000n V_low
+ 516.200001n V_low
+ 516.300000n V_low
+ 516.300001n V_low
+ 516.400000n V_low
+ 516.400001n V_low
+ 516.500000n V_low
+ 516.500001n V_low
+ 516.600000n V_low
+ 516.600001n V_low
+ 516.700000n V_low
+ 516.700001n V_low
+ 516.800000n V_low
+ 516.800001n V_low
+ 516.900000n V_low
+ 516.900001n V_low
+ 517.000000n V_low
+ 517.000001n V_low
+ 517.100000n V_low
+ 517.100001n V_low
+ 517.200000n V_low
+ 517.200001n V_low
+ 517.300000n V_low
+ 517.300001n V_low
+ 517.400000n V_low
+ 517.400001n V_low
+ 517.500000n V_low
+ 517.500001n V_low
+ 517.600000n V_low
+ 517.600001n V_low
+ 517.700000n V_low
+ 517.700001n V_low
+ 517.800000n V_low
+ 517.800001n V_low
+ 517.900000n V_low
+ 517.900001n V_low
+ 518.000000n V_low
+ 518.000001n V_low
+ 518.100000n V_low
+ 518.100001n V_low
+ 518.200000n V_low
+ 518.200001n V_low
+ 518.300000n V_low
+ 518.300001n V_low
+ 518.400000n V_low
+ 518.400001n V_low
+ 518.500000n V_low
+ 518.500001n V_low
+ 518.600000n V_low
+ 518.600001n V_low
+ 518.700000n V_low
+ 518.700001n V_low
+ 518.800000n V_low
+ 518.800001n V_low
+ 518.900000n V_low
+ 518.900001n V_low
+ 519.000000n V_low
+ 519.000001n V_low
+ 519.100000n V_low
+ 519.100001n V_low
+ 519.200000n V_low
+ 519.200001n V_low
+ 519.300000n V_low
+ 519.300001n V_low
+ 519.400000n V_low
+ 519.400001n V_low
+ 519.500000n V_low
+ 519.500001n V_low
+ 519.600000n V_low
+ 519.600001n V_low
+ 519.700000n V_low
+ 519.700001n V_low
+ 519.800000n V_low
+ 519.800001n V_low
+ 519.900000n V_low
+ 519.900001n V_low
+ 520.000000n V_low
+ 520.000001n V_hig
+ 520.100000n V_hig
+ 520.100001n V_hig
+ 520.200000n V_hig
+ 520.200001n V_hig
+ 520.300000n V_hig
+ 520.300001n V_hig
+ 520.400000n V_hig
+ 520.400001n V_hig
+ 520.500000n V_hig
+ 520.500001n V_hig
+ 520.600000n V_hig
+ 520.600001n V_hig
+ 520.700000n V_hig
+ 520.700001n V_hig
+ 520.800000n V_hig
+ 520.800001n V_hig
+ 520.900000n V_hig
+ 520.900001n V_hig
+ 521.000000n V_hig
+ 521.000001n V_low
+ 521.100000n V_low
+ 521.100001n V_low
+ 521.200000n V_low
+ 521.200001n V_low
+ 521.300000n V_low
+ 521.300001n V_low
+ 521.400000n V_low
+ 521.400001n V_low
+ 521.500000n V_low
+ 521.500001n V_low
+ 521.600000n V_low
+ 521.600001n V_low
+ 521.700000n V_low
+ 521.700001n V_low
+ 521.800000n V_low
+ 521.800001n V_low
+ 521.900000n V_low
+ 521.900001n V_low
+ 522.000000n V_low
+ 522.000001n V_hig
+ 522.100000n V_hig
+ 522.100001n V_hig
+ 522.200000n V_hig
+ 522.200001n V_hig
+ 522.300000n V_hig
+ 522.300001n V_hig
+ 522.400000n V_hig
+ 522.400001n V_hig
+ 522.500000n V_hig
+ 522.500001n V_hig
+ 522.600000n V_hig
+ 522.600001n V_hig
+ 522.700000n V_hig
+ 522.700001n V_hig
+ 522.800000n V_hig
+ 522.800001n V_hig
+ 522.900000n V_hig
+ 522.900001n V_hig
+ 523.000000n V_hig
+ 523.000001n V_hig
+ 523.100000n V_hig
+ 523.100001n V_hig
+ 523.200000n V_hig
+ 523.200001n V_hig
+ 523.300000n V_hig
+ 523.300001n V_hig
+ 523.400000n V_hig
+ 523.400001n V_hig
+ 523.500000n V_hig
+ 523.500001n V_hig
+ 523.600000n V_hig
+ 523.600001n V_hig
+ 523.700000n V_hig
+ 523.700001n V_hig
+ 523.800000n V_hig
+ 523.800001n V_hig
+ 523.900000n V_hig
+ 523.900001n V_hig
+ 524.000000n V_hig
+ 524.000001n V_low
+ 524.100000n V_low
+ 524.100001n V_low
+ 524.200000n V_low
+ 524.200001n V_low
+ 524.300000n V_low
+ 524.300001n V_low
+ 524.400000n V_low
+ 524.400001n V_low
+ 524.500000n V_low
+ 524.500001n V_low
+ 524.600000n V_low
+ 524.600001n V_low
+ 524.700000n V_low
+ 524.700001n V_low
+ 524.800000n V_low
+ 524.800001n V_low
+ 524.900000n V_low
+ 524.900001n V_low
+ 525.000000n V_low
+ 525.000001n V_hig
+ 525.100000n V_hig
+ 525.100001n V_hig
+ 525.200000n V_hig
+ 525.200001n V_hig
+ 525.300000n V_hig
+ 525.300001n V_hig
+ 525.400000n V_hig
+ 525.400001n V_hig
+ 525.500000n V_hig
+ 525.500001n V_hig
+ 525.600000n V_hig
+ 525.600001n V_hig
+ 525.700000n V_hig
+ 525.700001n V_hig
+ 525.800000n V_hig
+ 525.800001n V_hig
+ 525.900000n V_hig
+ 525.900001n V_hig
+ 526.000000n V_hig
+ 526.000001n V_low
+ 526.100000n V_low
+ 526.100001n V_low
+ 526.200000n V_low
+ 526.200001n V_low
+ 526.300000n V_low
+ 526.300001n V_low
+ 526.400000n V_low
+ 526.400001n V_low
+ 526.500000n V_low
+ 526.500001n V_low
+ 526.600000n V_low
+ 526.600001n V_low
+ 526.700000n V_low
+ 526.700001n V_low
+ 526.800000n V_low
+ 526.800001n V_low
+ 526.900000n V_low
+ 526.900001n V_low
+ 527.000000n V_low
+ 527.000001n V_hig
+ 527.100000n V_hig
+ 527.100001n V_hig
+ 527.200000n V_hig
+ 527.200001n V_hig
+ 527.300000n V_hig
+ 527.300001n V_hig
+ 527.400000n V_hig
+ 527.400001n V_hig
+ 527.500000n V_hig
+ 527.500001n V_hig
+ 527.600000n V_hig
+ 527.600001n V_hig
+ 527.700000n V_hig
+ 527.700001n V_hig
+ 527.800000n V_hig
+ 527.800001n V_hig
+ 527.900000n V_hig
+ 527.900001n V_hig
+ 528.000000n V_hig
+ 528.000001n V_low
+ 528.100000n V_low
+ 528.100001n V_low
+ 528.200000n V_low
+ 528.200001n V_low
+ 528.300000n V_low
+ 528.300001n V_low
+ 528.400000n V_low
+ 528.400001n V_low
+ 528.500000n V_low
+ 528.500001n V_low
+ 528.600000n V_low
+ 528.600001n V_low
+ 528.700000n V_low
+ 528.700001n V_low
+ 528.800000n V_low
+ 528.800001n V_low
+ 528.900000n V_low
+ 528.900001n V_low
+ 529.000000n V_low
+ 529.000001n V_hig
+ 529.100000n V_hig
+ 529.100001n V_hig
+ 529.200000n V_hig
+ 529.200001n V_hig
+ 529.300000n V_hig
+ 529.300001n V_hig
+ 529.400000n V_hig
+ 529.400001n V_hig
+ 529.500000n V_hig
+ 529.500001n V_hig
+ 529.600000n V_hig
+ 529.600001n V_hig
+ 529.700000n V_hig
+ 529.700001n V_hig
+ 529.800000n V_hig
+ 529.800001n V_hig
+ 529.900000n V_hig
+ 529.900001n V_hig
+ 530.000000n V_hig
+ 530.000001n V_low
+ 530.100000n V_low
+ 530.100001n V_low
+ 530.200000n V_low
+ 530.200001n V_low
+ 530.300000n V_low
+ 530.300001n V_low
+ 530.400000n V_low
+ 530.400001n V_low
+ 530.500000n V_low
+ 530.500001n V_low
+ 530.600000n V_low
+ 530.600001n V_low
+ 530.700000n V_low
+ 530.700001n V_low
+ 530.800000n V_low
+ 530.800001n V_low
+ 530.900000n V_low
+ 530.900001n V_low
+ 531.000000n V_low
+ 531.000001n V_low
+ 531.100000n V_low
+ 531.100001n V_low
+ 531.200000n V_low
+ 531.200001n V_low
+ 531.300000n V_low
+ 531.300001n V_low
+ 531.400000n V_low
+ 531.400001n V_low
+ 531.500000n V_low
+ 531.500001n V_low
+ 531.600000n V_low
+ 531.600001n V_low
+ 531.700000n V_low
+ 531.700001n V_low
+ 531.800000n V_low
+ 531.800001n V_low
+ 531.900000n V_low
+ 531.900001n V_low
+ 532.000000n V_low
+ 532.000001n V_hig
+ 532.100000n V_hig
+ 532.100001n V_hig
+ 532.200000n V_hig
+ 532.200001n V_hig
+ 532.300000n V_hig
+ 532.300001n V_hig
+ 532.400000n V_hig
+ 532.400001n V_hig
+ 532.500000n V_hig
+ 532.500001n V_hig
+ 532.600000n V_hig
+ 532.600001n V_hig
+ 532.700000n V_hig
+ 532.700001n V_hig
+ 532.800000n V_hig
+ 532.800001n V_hig
+ 532.900000n V_hig
+ 532.900001n V_hig
+ 533.000000n V_hig
+ 533.000001n V_hig
+ 533.100000n V_hig
+ 533.100001n V_hig
+ 533.200000n V_hig
+ 533.200001n V_hig
+ 533.300000n V_hig
+ 533.300001n V_hig
+ 533.400000n V_hig
+ 533.400001n V_hig
+ 533.500000n V_hig
+ 533.500001n V_hig
+ 533.600000n V_hig
+ 533.600001n V_hig
+ 533.700000n V_hig
+ 533.700001n V_hig
+ 533.800000n V_hig
+ 533.800001n V_hig
+ 533.900000n V_hig
+ 533.900001n V_hig
+ 534.000000n V_hig
+ 534.000001n V_hig
+ 534.100000n V_hig
+ 534.100001n V_hig
+ 534.200000n V_hig
+ 534.200001n V_hig
+ 534.300000n V_hig
+ 534.300001n V_hig
+ 534.400000n V_hig
+ 534.400001n V_hig
+ 534.500000n V_hig
+ 534.500001n V_hig
+ 534.600000n V_hig
+ 534.600001n V_hig
+ 534.700000n V_hig
+ 534.700001n V_hig
+ 534.800000n V_hig
+ 534.800001n V_hig
+ 534.900000n V_hig
+ 534.900001n V_hig
+ 535.000000n V_hig
+ 535.000001n V_hig
+ 535.100000n V_hig
+ 535.100001n V_hig
+ 535.200000n V_hig
+ 535.200001n V_hig
+ 535.300000n V_hig
+ 535.300001n V_hig
+ 535.400000n V_hig
+ 535.400001n V_hig
+ 535.500000n V_hig
+ 535.500001n V_hig
+ 535.600000n V_hig
+ 535.600001n V_hig
+ 535.700000n V_hig
+ 535.700001n V_hig
+ 535.800000n V_hig
+ 535.800001n V_hig
+ 535.900000n V_hig
+ 535.900001n V_hig
+ 536.000000n V_hig
+ 536.000001n V_hig
+ 536.100000n V_hig
+ 536.100001n V_hig
+ 536.200000n V_hig
+ 536.200001n V_hig
+ 536.300000n V_hig
+ 536.300001n V_hig
+ 536.400000n V_hig
+ 536.400001n V_hig
+ 536.500000n V_hig
+ 536.500001n V_hig
+ 536.600000n V_hig
+ 536.600001n V_hig
+ 536.700000n V_hig
+ 536.700001n V_hig
+ 536.800000n V_hig
+ 536.800001n V_hig
+ 536.900000n V_hig
+ 536.900001n V_hig
+ 537.000000n V_hig
+ 537.000001n V_hig
+ 537.100000n V_hig
+ 537.100001n V_hig
+ 537.200000n V_hig
+ 537.200001n V_hig
+ 537.300000n V_hig
+ 537.300001n V_hig
+ 537.400000n V_hig
+ 537.400001n V_hig
+ 537.500000n V_hig
+ 537.500001n V_hig
+ 537.600000n V_hig
+ 537.600001n V_hig
+ 537.700000n V_hig
+ 537.700001n V_hig
+ 537.800000n V_hig
+ 537.800001n V_hig
+ 537.900000n V_hig
+ 537.900001n V_hig
+ 538.000000n V_hig
+ 538.000001n V_low
+ 538.100000n V_low
+ 538.100001n V_low
+ 538.200000n V_low
+ 538.200001n V_low
+ 538.300000n V_low
+ 538.300001n V_low
+ 538.400000n V_low
+ 538.400001n V_low
+ 538.500000n V_low
+ 538.500001n V_low
+ 538.600000n V_low
+ 538.600001n V_low
+ 538.700000n V_low
+ 538.700001n V_low
+ 538.800000n V_low
+ 538.800001n V_low
+ 538.900000n V_low
+ 538.900001n V_low
+ 539.000000n V_low
+ 539.000001n V_hig
+ 539.100000n V_hig
+ 539.100001n V_hig
+ 539.200000n V_hig
+ 539.200001n V_hig
+ 539.300000n V_hig
+ 539.300001n V_hig
+ 539.400000n V_hig
+ 539.400001n V_hig
+ 539.500000n V_hig
+ 539.500001n V_hig
+ 539.600000n V_hig
+ 539.600001n V_hig
+ 539.700000n V_hig
+ 539.700001n V_hig
+ 539.800000n V_hig
+ 539.800001n V_hig
+ 539.900000n V_hig
+ 539.900001n V_hig
+ 540.000000n V_hig
+ 540.000001n V_low
+ 540.100000n V_low
+ 540.100001n V_low
+ 540.200000n V_low
+ 540.200001n V_low
+ 540.300000n V_low
+ 540.300001n V_low
+ 540.400000n V_low
+ 540.400001n V_low
+ 540.500000n V_low
+ 540.500001n V_low
+ 540.600000n V_low
+ 540.600001n V_low
+ 540.700000n V_low
+ 540.700001n V_low
+ 540.800000n V_low
+ 540.800001n V_low
+ 540.900000n V_low
+ 540.900001n V_low
+ 541.000000n V_low
+ 541.000001n V_low
+ 541.100000n V_low
+ 541.100001n V_low
+ 541.200000n V_low
+ 541.200001n V_low
+ 541.300000n V_low
+ 541.300001n V_low
+ 541.400000n V_low
+ 541.400001n V_low
+ 541.500000n V_low
+ 541.500001n V_low
+ 541.600000n V_low
+ 541.600001n V_low
+ 541.700000n V_low
+ 541.700001n V_low
+ 541.800000n V_low
+ 541.800001n V_low
+ 541.900000n V_low
+ 541.900001n V_low
+ 542.000000n V_low
+ 542.000001n V_low
+ 542.100000n V_low
+ 542.100001n V_low
+ 542.200000n V_low
+ 542.200001n V_low
+ 542.300000n V_low
+ 542.300001n V_low
+ 542.400000n V_low
+ 542.400001n V_low
+ 542.500000n V_low
+ 542.500001n V_low
+ 542.600000n V_low
+ 542.600001n V_low
+ 542.700000n V_low
+ 542.700001n V_low
+ 542.800000n V_low
+ 542.800001n V_low
+ 542.900000n V_low
+ 542.900001n V_low
+ 543.000000n V_low
+ 543.000001n V_hig
+ 543.100000n V_hig
+ 543.100001n V_hig
+ 543.200000n V_hig
+ 543.200001n V_hig
+ 543.300000n V_hig
+ 543.300001n V_hig
+ 543.400000n V_hig
+ 543.400001n V_hig
+ 543.500000n V_hig
+ 543.500001n V_hig
+ 543.600000n V_hig
+ 543.600001n V_hig
+ 543.700000n V_hig
+ 543.700001n V_hig
+ 543.800000n V_hig
+ 543.800001n V_hig
+ 543.900000n V_hig
+ 543.900001n V_hig
+ 544.000000n V_hig
+ 544.000001n V_low
+ 544.100000n V_low
+ 544.100001n V_low
+ 544.200000n V_low
+ 544.200001n V_low
+ 544.300000n V_low
+ 544.300001n V_low
+ 544.400000n V_low
+ 544.400001n V_low
+ 544.500000n V_low
+ 544.500001n V_low
+ 544.600000n V_low
+ 544.600001n V_low
+ 544.700000n V_low
+ 544.700001n V_low
+ 544.800000n V_low
+ 544.800001n V_low
+ 544.900000n V_low
+ 544.900001n V_low
+ 545.000000n V_low
+ 545.000001n V_low
+ 545.100000n V_low
+ 545.100001n V_low
+ 545.200000n V_low
+ 545.200001n V_low
+ 545.300000n V_low
+ 545.300001n V_low
+ 545.400000n V_low
+ 545.400001n V_low
+ 545.500000n V_low
+ 545.500001n V_low
+ 545.600000n V_low
+ 545.600001n V_low
+ 545.700000n V_low
+ 545.700001n V_low
+ 545.800000n V_low
+ 545.800001n V_low
+ 545.900000n V_low
+ 545.900001n V_low
+ 546.000000n V_low
+ 546.000001n V_hig
+ 546.100000n V_hig
+ 546.100001n V_hig
+ 546.200000n V_hig
+ 546.200001n V_hig
+ 546.300000n V_hig
+ 546.300001n V_hig
+ 546.400000n V_hig
+ 546.400001n V_hig
+ 546.500000n V_hig
+ 546.500001n V_hig
+ 546.600000n V_hig
+ 546.600001n V_hig
+ 546.700000n V_hig
+ 546.700001n V_hig
+ 546.800000n V_hig
+ 546.800001n V_hig
+ 546.900000n V_hig
+ 546.900001n V_hig
+ 547.000000n V_hig
+ 547.000001n V_hig
+ 547.100000n V_hig
+ 547.100001n V_hig
+ 547.200000n V_hig
+ 547.200001n V_hig
+ 547.300000n V_hig
+ 547.300001n V_hig
+ 547.400000n V_hig
+ 547.400001n V_hig
+ 547.500000n V_hig
+ 547.500001n V_hig
+ 547.600000n V_hig
+ 547.600001n V_hig
+ 547.700000n V_hig
+ 547.700001n V_hig
+ 547.800000n V_hig
+ 547.800001n V_hig
+ 547.900000n V_hig
+ 547.900001n V_hig
+ 548.000000n V_hig
+ 548.000001n V_low
+ 548.100000n V_low
+ 548.100001n V_low
+ 548.200000n V_low
+ 548.200001n V_low
+ 548.300000n V_low
+ 548.300001n V_low
+ 548.400000n V_low
+ 548.400001n V_low
+ 548.500000n V_low
+ 548.500001n V_low
+ 548.600000n V_low
+ 548.600001n V_low
+ 548.700000n V_low
+ 548.700001n V_low
+ 548.800000n V_low
+ 548.800001n V_low
+ 548.900000n V_low
+ 548.900001n V_low
+ 549.000000n V_low
+ 549.000001n V_hig
+ 549.100000n V_hig
+ 549.100001n V_hig
+ 549.200000n V_hig
+ 549.200001n V_hig
+ 549.300000n V_hig
+ 549.300001n V_hig
+ 549.400000n V_hig
+ 549.400001n V_hig
+ 549.500000n V_hig
+ 549.500001n V_hig
+ 549.600000n V_hig
+ 549.600001n V_hig
+ 549.700000n V_hig
+ 549.700001n V_hig
+ 549.800000n V_hig
+ 549.800001n V_hig
+ 549.900000n V_hig
+ 549.900001n V_hig
+ 550.000000n V_hig
+ 550.000001n V_hig
+ 550.100000n V_hig
+ 550.100001n V_hig
+ 550.200000n V_hig
+ 550.200001n V_hig
+ 550.300000n V_hig
+ 550.300001n V_hig
+ 550.400000n V_hig
+ 550.400001n V_hig
+ 550.500000n V_hig
+ 550.500001n V_hig
+ 550.600000n V_hig
+ 550.600001n V_hig
+ 550.700000n V_hig
+ 550.700001n V_hig
+ 550.800000n V_hig
+ 550.800001n V_hig
+ 550.900000n V_hig
+ 550.900001n V_hig
+ 551.000000n V_hig
+ 551.000001n V_low
+ 551.100000n V_low
+ 551.100001n V_low
+ 551.200000n V_low
+ 551.200001n V_low
+ 551.300000n V_low
+ 551.300001n V_low
+ 551.400000n V_low
+ 551.400001n V_low
+ 551.500000n V_low
+ 551.500001n V_low
+ 551.600000n V_low
+ 551.600001n V_low
+ 551.700000n V_low
+ 551.700001n V_low
+ 551.800000n V_low
+ 551.800001n V_low
+ 551.900000n V_low
+ 551.900001n V_low
+ 552.000000n V_low
+ 552.000001n V_low
+ 552.100000n V_low
+ 552.100001n V_low
+ 552.200000n V_low
+ 552.200001n V_low
+ 552.300000n V_low
+ 552.300001n V_low
+ 552.400000n V_low
+ 552.400001n V_low
+ 552.500000n V_low
+ 552.500001n V_low
+ 552.600000n V_low
+ 552.600001n V_low
+ 552.700000n V_low
+ 552.700001n V_low
+ 552.800000n V_low
+ 552.800001n V_low
+ 552.900000n V_low
+ 552.900001n V_low
+ 553.000000n V_low
+ 553.000001n V_low
+ 553.100000n V_low
+ 553.100001n V_low
+ 553.200000n V_low
+ 553.200001n V_low
+ 553.300000n V_low
+ 553.300001n V_low
+ 553.400000n V_low
+ 553.400001n V_low
+ 553.500000n V_low
+ 553.500001n V_low
+ 553.600000n V_low
+ 553.600001n V_low
+ 553.700000n V_low
+ 553.700001n V_low
+ 553.800000n V_low
+ 553.800001n V_low
+ 553.900000n V_low
+ 553.900001n V_low
+ 554.000000n V_low
+ 554.000001n V_hig
+ 554.100000n V_hig
+ 554.100001n V_hig
+ 554.200000n V_hig
+ 554.200001n V_hig
+ 554.300000n V_hig
+ 554.300001n V_hig
+ 554.400000n V_hig
+ 554.400001n V_hig
+ 554.500000n V_hig
+ 554.500001n V_hig
+ 554.600000n V_hig
+ 554.600001n V_hig
+ 554.700000n V_hig
+ 554.700001n V_hig
+ 554.800000n V_hig
+ 554.800001n V_hig
+ 554.900000n V_hig
+ 554.900001n V_hig
+ 555.000000n V_hig
+ 555.000001n V_low
+ 555.100000n V_low
+ 555.100001n V_low
+ 555.200000n V_low
+ 555.200001n V_low
+ 555.300000n V_low
+ 555.300001n V_low
+ 555.400000n V_low
+ 555.400001n V_low
+ 555.500000n V_low
+ 555.500001n V_low
+ 555.600000n V_low
+ 555.600001n V_low
+ 555.700000n V_low
+ 555.700001n V_low
+ 555.800000n V_low
+ 555.800001n V_low
+ 555.900000n V_low
+ 555.900001n V_low
+ 556.000000n V_low
+ 556.000001n V_hig
+ 556.100000n V_hig
+ 556.100001n V_hig
+ 556.200000n V_hig
+ 556.200001n V_hig
+ 556.300000n V_hig
+ 556.300001n V_hig
+ 556.400000n V_hig
+ 556.400001n V_hig
+ 556.500000n V_hig
+ 556.500001n V_hig
+ 556.600000n V_hig
+ 556.600001n V_hig
+ 556.700000n V_hig
+ 556.700001n V_hig
+ 556.800000n V_hig
+ 556.800001n V_hig
+ 556.900000n V_hig
+ 556.900001n V_hig
+ 557.000000n V_hig
+ 557.000001n V_low
+ 557.100000n V_low
+ 557.100001n V_low
+ 557.200000n V_low
+ 557.200001n V_low
+ 557.300000n V_low
+ 557.300001n V_low
+ 557.400000n V_low
+ 557.400001n V_low
+ 557.500000n V_low
+ 557.500001n V_low
+ 557.600000n V_low
+ 557.600001n V_low
+ 557.700000n V_low
+ 557.700001n V_low
+ 557.800000n V_low
+ 557.800001n V_low
+ 557.900000n V_low
+ 557.900001n V_low
+ 558.000000n V_low
+ 558.000001n V_low
+ 558.100000n V_low
+ 558.100001n V_low
+ 558.200000n V_low
+ 558.200001n V_low
+ 558.300000n V_low
+ 558.300001n V_low
+ 558.400000n V_low
+ 558.400001n V_low
+ 558.500000n V_low
+ 558.500001n V_low
+ 558.600000n V_low
+ 558.600001n V_low
+ 558.700000n V_low
+ 558.700001n V_low
+ 558.800000n V_low
+ 558.800001n V_low
+ 558.900000n V_low
+ 558.900001n V_low
+ 559.000000n V_low
+ 559.000001n V_low
+ 559.100000n V_low
+ 559.100001n V_low
+ 559.200000n V_low
+ 559.200001n V_low
+ 559.300000n V_low
+ 559.300001n V_low
+ 559.400000n V_low
+ 559.400001n V_low
+ 559.500000n V_low
+ 559.500001n V_low
+ 559.600000n V_low
+ 559.600001n V_low
+ 559.700000n V_low
+ 559.700001n V_low
+ 559.800000n V_low
+ 559.800001n V_low
+ 559.900000n V_low
+ 559.900001n V_low
+ 560.000000n V_low
+ 560.000001n V_low
+ 560.100000n V_low
+ 560.100001n V_low
+ 560.200000n V_low
+ 560.200001n V_low
+ 560.300000n V_low
+ 560.300001n V_low
+ 560.400000n V_low
+ 560.400001n V_low
+ 560.500000n V_low
+ 560.500001n V_low
+ 560.600000n V_low
+ 560.600001n V_low
+ 560.700000n V_low
+ 560.700001n V_low
+ 560.800000n V_low
+ 560.800001n V_low
+ 560.900000n V_low
+ 560.900001n V_low
+ 561.000000n V_low
+ 561.000001n V_low
+ 561.100000n V_low
+ 561.100001n V_low
+ 561.200000n V_low
+ 561.200001n V_low
+ 561.300000n V_low
+ 561.300001n V_low
+ 561.400000n V_low
+ 561.400001n V_low
+ 561.500000n V_low
+ 561.500001n V_low
+ 561.600000n V_low
+ 561.600001n V_low
+ 561.700000n V_low
+ 561.700001n V_low
+ 561.800000n V_low
+ 561.800001n V_low
+ 561.900000n V_low
+ 561.900001n V_low
+ 562.000000n V_low
+ 562.000001n V_low
+ 562.100000n V_low
+ 562.100001n V_low
+ 562.200000n V_low
+ 562.200001n V_low
+ 562.300000n V_low
+ 562.300001n V_low
+ 562.400000n V_low
+ 562.400001n V_low
+ 562.500000n V_low
+ 562.500001n V_low
+ 562.600000n V_low
+ 562.600001n V_low
+ 562.700000n V_low
+ 562.700001n V_low
+ 562.800000n V_low
+ 562.800001n V_low
+ 562.900000n V_low
+ 562.900001n V_low
+ 563.000000n V_low
+ 563.000001n V_hig
+ 563.100000n V_hig
+ 563.100001n V_hig
+ 563.200000n V_hig
+ 563.200001n V_hig
+ 563.300000n V_hig
+ 563.300001n V_hig
+ 563.400000n V_hig
+ 563.400001n V_hig
+ 563.500000n V_hig
+ 563.500001n V_hig
+ 563.600000n V_hig
+ 563.600001n V_hig
+ 563.700000n V_hig
+ 563.700001n V_hig
+ 563.800000n V_hig
+ 563.800001n V_hig
+ 563.900000n V_hig
+ 563.900001n V_hig
+ 564.000000n V_hig
+ 564.000001n V_low
+ 564.100000n V_low
+ 564.100001n V_low
+ 564.200000n V_low
+ 564.200001n V_low
+ 564.300000n V_low
+ 564.300001n V_low
+ 564.400000n V_low
+ 564.400001n V_low
+ 564.500000n V_low
+ 564.500001n V_low
+ 564.600000n V_low
+ 564.600001n V_low
+ 564.700000n V_low
+ 564.700001n V_low
+ 564.800000n V_low
+ 564.800001n V_low
+ 564.900000n V_low
+ 564.900001n V_low
+ 565.000000n V_low
+ 565.000001n V_low
+ 565.100000n V_low
+ 565.100001n V_low
+ 565.200000n V_low
+ 565.200001n V_low
+ 565.300000n V_low
+ 565.300001n V_low
+ 565.400000n V_low
+ 565.400001n V_low
+ 565.500000n V_low
+ 565.500001n V_low
+ 565.600000n V_low
+ 565.600001n V_low
+ 565.700000n V_low
+ 565.700001n V_low
+ 565.800000n V_low
+ 565.800001n V_low
+ 565.900000n V_low
+ 565.900001n V_low
+ 566.000000n V_low
+ 566.000001n V_low
+ 566.100000n V_low
+ 566.100001n V_low
+ 566.200000n V_low
+ 566.200001n V_low
+ 566.300000n V_low
+ 566.300001n V_low
+ 566.400000n V_low
+ 566.400001n V_low
+ 566.500000n V_low
+ 566.500001n V_low
+ 566.600000n V_low
+ 566.600001n V_low
+ 566.700000n V_low
+ 566.700001n V_low
+ 566.800000n V_low
+ 566.800001n V_low
+ 566.900000n V_low
+ 566.900001n V_low
+ 567.000000n V_low
+ 567.000001n V_low
+ 567.100000n V_low
+ 567.100001n V_low
+ 567.200000n V_low
+ 567.200001n V_low
+ 567.300000n V_low
+ 567.300001n V_low
+ 567.400000n V_low
+ 567.400001n V_low
+ 567.500000n V_low
+ 567.500001n V_low
+ 567.600000n V_low
+ 567.600001n V_low
+ 567.700000n V_low
+ 567.700001n V_low
+ 567.800000n V_low
+ 567.800001n V_low
+ 567.900000n V_low
+ 567.900001n V_low
+ 568.000000n V_low
+ 568.000001n V_low
+ 568.100000n V_low
+ 568.100001n V_low
+ 568.200000n V_low
+ 568.200001n V_low
+ 568.300000n V_low
+ 568.300001n V_low
+ 568.400000n V_low
+ 568.400001n V_low
+ 568.500000n V_low
+ 568.500001n V_low
+ 568.600000n V_low
+ 568.600001n V_low
+ 568.700000n V_low
+ 568.700001n V_low
+ 568.800000n V_low
+ 568.800001n V_low
+ 568.900000n V_low
+ 568.900001n V_low
+ 569.000000n V_low
+ 569.000001n V_hig
+ 569.100000n V_hig
+ 569.100001n V_hig
+ 569.200000n V_hig
+ 569.200001n V_hig
+ 569.300000n V_hig
+ 569.300001n V_hig
+ 569.400000n V_hig
+ 569.400001n V_hig
+ 569.500000n V_hig
+ 569.500001n V_hig
+ 569.600000n V_hig
+ 569.600001n V_hig
+ 569.700000n V_hig
+ 569.700001n V_hig
+ 569.800000n V_hig
+ 569.800001n V_hig
+ 569.900000n V_hig
+ 569.900001n V_hig
+ 570.000000n V_hig
+ 570.000001n V_hig
+ 570.100000n V_hig
+ 570.100001n V_hig
+ 570.200000n V_hig
+ 570.200001n V_hig
+ 570.300000n V_hig
+ 570.300001n V_hig
+ 570.400000n V_hig
+ 570.400001n V_hig
+ 570.500000n V_hig
+ 570.500001n V_hig
+ 570.600000n V_hig
+ 570.600001n V_hig
+ 570.700000n V_hig
+ 570.700001n V_hig
+ 570.800000n V_hig
+ 570.800001n V_hig
+ 570.900000n V_hig
+ 570.900001n V_hig
+ 571.000000n V_hig
+ 571.000001n V_hig
+ 571.100000n V_hig
+ 571.100001n V_hig
+ 571.200000n V_hig
+ 571.200001n V_hig
+ 571.300000n V_hig
+ 571.300001n V_hig
+ 571.400000n V_hig
+ 571.400001n V_hig
+ 571.500000n V_hig
+ 571.500001n V_hig
+ 571.600000n V_hig
+ 571.600001n V_hig
+ 571.700000n V_hig
+ 571.700001n V_hig
+ 571.800000n V_hig
+ 571.800001n V_hig
+ 571.900000n V_hig
+ 571.900001n V_hig
+ 572.000000n V_hig
+ 572.000001n V_hig
+ 572.100000n V_hig
+ 572.100001n V_hig
+ 572.200000n V_hig
+ 572.200001n V_hig
+ 572.300000n V_hig
+ 572.300001n V_hig
+ 572.400000n V_hig
+ 572.400001n V_hig
+ 572.500000n V_hig
+ 572.500001n V_hig
+ 572.600000n V_hig
+ 572.600001n V_hig
+ 572.700000n V_hig
+ 572.700001n V_hig
+ 572.800000n V_hig
+ 572.800001n V_hig
+ 572.900000n V_hig
+ 572.900001n V_hig
+ 573.000000n V_hig
+ 573.000001n V_hig
+ 573.100000n V_hig
+ 573.100001n V_hig
+ 573.200000n V_hig
+ 573.200001n V_hig
+ 573.300000n V_hig
+ 573.300001n V_hig
+ 573.400000n V_hig
+ 573.400001n V_hig
+ 573.500000n V_hig
+ 573.500001n V_hig
+ 573.600000n V_hig
+ 573.600001n V_hig
+ 573.700000n V_hig
+ 573.700001n V_hig
+ 573.800000n V_hig
+ 573.800001n V_hig
+ 573.900000n V_hig
+ 573.900001n V_hig
+ 574.000000n V_hig
+ 574.000001n V_low
+ 574.100000n V_low
+ 574.100001n V_low
+ 574.200000n V_low
+ 574.200001n V_low
+ 574.300000n V_low
+ 574.300001n V_low
+ 574.400000n V_low
+ 574.400001n V_low
+ 574.500000n V_low
+ 574.500001n V_low
+ 574.600000n V_low
+ 574.600001n V_low
+ 574.700000n V_low
+ 574.700001n V_low
+ 574.800000n V_low
+ 574.800001n V_low
+ 574.900000n V_low
+ 574.900001n V_low
+ 575.000000n V_low
+ 575.000001n V_low
+ 575.100000n V_low
+ 575.100001n V_low
+ 575.200000n V_low
+ 575.200001n V_low
+ 575.300000n V_low
+ 575.300001n V_low
+ 575.400000n V_low
+ 575.400001n V_low
+ 575.500000n V_low
+ 575.500001n V_low
+ 575.600000n V_low
+ 575.600001n V_low
+ 575.700000n V_low
+ 575.700001n V_low
+ 575.800000n V_low
+ 575.800001n V_low
+ 575.900000n V_low
+ 575.900001n V_low
+ 576.000000n V_low
+ 576.000001n V_hig
+ 576.100000n V_hig
+ 576.100001n V_hig
+ 576.200000n V_hig
+ 576.200001n V_hig
+ 576.300000n V_hig
+ 576.300001n V_hig
+ 576.400000n V_hig
+ 576.400001n V_hig
+ 576.500000n V_hig
+ 576.500001n V_hig
+ 576.600000n V_hig
+ 576.600001n V_hig
+ 576.700000n V_hig
+ 576.700001n V_hig
+ 576.800000n V_hig
+ 576.800001n V_hig
+ 576.900000n V_hig
+ 576.900001n V_hig
+ 577.000000n V_hig
+ 577.000001n V_hig
+ 577.100000n V_hig
+ 577.100001n V_hig
+ 577.200000n V_hig
+ 577.200001n V_hig
+ 577.300000n V_hig
+ 577.300001n V_hig
+ 577.400000n V_hig
+ 577.400001n V_hig
+ 577.500000n V_hig
+ 577.500001n V_hig
+ 577.600000n V_hig
+ 577.600001n V_hig
+ 577.700000n V_hig
+ 577.700001n V_hig
+ 577.800000n V_hig
+ 577.800001n V_hig
+ 577.900000n V_hig
+ 577.900001n V_hig
+ 578.000000n V_hig
+ 578.000001n V_low
+ 578.100000n V_low
+ 578.100001n V_low
+ 578.200000n V_low
+ 578.200001n V_low
+ 578.300000n V_low
+ 578.300001n V_low
+ 578.400000n V_low
+ 578.400001n V_low
+ 578.500000n V_low
+ 578.500001n V_low
+ 578.600000n V_low
+ 578.600001n V_low
+ 578.700000n V_low
+ 578.700001n V_low
+ 578.800000n V_low
+ 578.800001n V_low
+ 578.900000n V_low
+ 578.900001n V_low
+ 579.000000n V_low
+ 579.000001n V_hig
+ 579.100000n V_hig
+ 579.100001n V_hig
+ 579.200000n V_hig
+ 579.200001n V_hig
+ 579.300000n V_hig
+ 579.300001n V_hig
+ 579.400000n V_hig
+ 579.400001n V_hig
+ 579.500000n V_hig
+ 579.500001n V_hig
+ 579.600000n V_hig
+ 579.600001n V_hig
+ 579.700000n V_hig
+ 579.700001n V_hig
+ 579.800000n V_hig
+ 579.800001n V_hig
+ 579.900000n V_hig
+ 579.900001n V_hig
+ 580.000000n V_hig
+ 580.000001n V_low
+ 580.100000n V_low
+ 580.100001n V_low
+ 580.200000n V_low
+ 580.200001n V_low
+ 580.300000n V_low
+ 580.300001n V_low
+ 580.400000n V_low
+ 580.400001n V_low
+ 580.500000n V_low
+ 580.500001n V_low
+ 580.600000n V_low
+ 580.600001n V_low
+ 580.700000n V_low
+ 580.700001n V_low
+ 580.800000n V_low
+ 580.800001n V_low
+ 580.900000n V_low
+ 580.900001n V_low
+ 581.000000n V_low
+ 581.000001n V_low
+ 581.100000n V_low
+ 581.100001n V_low
+ 581.200000n V_low
+ 581.200001n V_low
+ 581.300000n V_low
+ 581.300001n V_low
+ 581.400000n V_low
+ 581.400001n V_low
+ 581.500000n V_low
+ 581.500001n V_low
+ 581.600000n V_low
+ 581.600001n V_low
+ 581.700000n V_low
+ 581.700001n V_low
+ 581.800000n V_low
+ 581.800001n V_low
+ 581.900000n V_low
+ 581.900001n V_low
+ 582.000000n V_low
+ 582.000001n V_hig
+ 582.100000n V_hig
+ 582.100001n V_hig
+ 582.200000n V_hig
+ 582.200001n V_hig
+ 582.300000n V_hig
+ 582.300001n V_hig
+ 582.400000n V_hig
+ 582.400001n V_hig
+ 582.500000n V_hig
+ 582.500001n V_hig
+ 582.600000n V_hig
+ 582.600001n V_hig
+ 582.700000n V_hig
+ 582.700001n V_hig
+ 582.800000n V_hig
+ 582.800001n V_hig
+ 582.900000n V_hig
+ 582.900001n V_hig
+ 583.000000n V_hig
+ 583.000001n V_hig
+ 583.100000n V_hig
+ 583.100001n V_hig
+ 583.200000n V_hig
+ 583.200001n V_hig
+ 583.300000n V_hig
+ 583.300001n V_hig
+ 583.400000n V_hig
+ 583.400001n V_hig
+ 583.500000n V_hig
+ 583.500001n V_hig
+ 583.600000n V_hig
+ 583.600001n V_hig
+ 583.700000n V_hig
+ 583.700001n V_hig
+ 583.800000n V_hig
+ 583.800001n V_hig
+ 583.900000n V_hig
+ 583.900001n V_hig
+ 584.000000n V_hig
+ 584.000001n V_hig
+ 584.100000n V_hig
+ 584.100001n V_hig
+ 584.200000n V_hig
+ 584.200001n V_hig
+ 584.300000n V_hig
+ 584.300001n V_hig
+ 584.400000n V_hig
+ 584.400001n V_hig
+ 584.500000n V_hig
+ 584.500001n V_hig
+ 584.600000n V_hig
+ 584.600001n V_hig
+ 584.700000n V_hig
+ 584.700001n V_hig
+ 584.800000n V_hig
+ 584.800001n V_hig
+ 584.900000n V_hig
+ 584.900001n V_hig
+ 585.000000n V_hig
+ 585.000001n V_hig
+ 585.100000n V_hig
+ 585.100001n V_hig
+ 585.200000n V_hig
+ 585.200001n V_hig
+ 585.300000n V_hig
+ 585.300001n V_hig
+ 585.400000n V_hig
+ 585.400001n V_hig
+ 585.500000n V_hig
+ 585.500001n V_hig
+ 585.600000n V_hig
+ 585.600001n V_hig
+ 585.700000n V_hig
+ 585.700001n V_hig
+ 585.800000n V_hig
+ 585.800001n V_hig
+ 585.900000n V_hig
+ 585.900001n V_hig
+ 586.000000n V_hig
+ 586.000001n V_hig
+ 586.100000n V_hig
+ 586.100001n V_hig
+ 586.200000n V_hig
+ 586.200001n V_hig
+ 586.300000n V_hig
+ 586.300001n V_hig
+ 586.400000n V_hig
+ 586.400001n V_hig
+ 586.500000n V_hig
+ 586.500001n V_hig
+ 586.600000n V_hig
+ 586.600001n V_hig
+ 586.700000n V_hig
+ 586.700001n V_hig
+ 586.800000n V_hig
+ 586.800001n V_hig
+ 586.900000n V_hig
+ 586.900001n V_hig
+ 587.000000n V_hig
+ 587.000001n V_low
+ 587.100000n V_low
+ 587.100001n V_low
+ 587.200000n V_low
+ 587.200001n V_low
+ 587.300000n V_low
+ 587.300001n V_low
+ 587.400000n V_low
+ 587.400001n V_low
+ 587.500000n V_low
+ 587.500001n V_low
+ 587.600000n V_low
+ 587.600001n V_low
+ 587.700000n V_low
+ 587.700001n V_low
+ 587.800000n V_low
+ 587.800001n V_low
+ 587.900000n V_low
+ 587.900001n V_low
+ 588.000000n V_low
+ 588.000001n V_hig
+ 588.100000n V_hig
+ 588.100001n V_hig
+ 588.200000n V_hig
+ 588.200001n V_hig
+ 588.300000n V_hig
+ 588.300001n V_hig
+ 588.400000n V_hig
+ 588.400001n V_hig
+ 588.500000n V_hig
+ 588.500001n V_hig
+ 588.600000n V_hig
+ 588.600001n V_hig
+ 588.700000n V_hig
+ 588.700001n V_hig
+ 588.800000n V_hig
+ 588.800001n V_hig
+ 588.900000n V_hig
+ 588.900001n V_hig
+ 589.000000n V_hig
+ 589.000001n V_low
+ 589.100000n V_low
+ 589.100001n V_low
+ 589.200000n V_low
+ 589.200001n V_low
+ 589.300000n V_low
+ 589.300001n V_low
+ 589.400000n V_low
+ 589.400001n V_low
+ 589.500000n V_low
+ 589.500001n V_low
+ 589.600000n V_low
+ 589.600001n V_low
+ 589.700000n V_low
+ 589.700001n V_low
+ 589.800000n V_low
+ 589.800001n V_low
+ 589.900000n V_low
+ 589.900001n V_low
+ 590.000000n V_low
+ 590.000001n V_low
+ 590.100000n V_low
+ 590.100001n V_low
+ 590.200000n V_low
+ 590.200001n V_low
+ 590.300000n V_low
+ 590.300001n V_low
+ 590.400000n V_low
+ 590.400001n V_low
+ 590.500000n V_low
+ 590.500001n V_low
+ 590.600000n V_low
+ 590.600001n V_low
+ 590.700000n V_low
+ 590.700001n V_low
+ 590.800000n V_low
+ 590.800001n V_low
+ 590.900000n V_low
+ 590.900001n V_low
+ 591.000000n V_low
+ 591.000001n V_low
+ 591.100000n V_low
+ 591.100001n V_low
+ 591.200000n V_low
+ 591.200001n V_low
+ 591.300000n V_low
+ 591.300001n V_low
+ 591.400000n V_low
+ 591.400001n V_low
+ 591.500000n V_low
+ 591.500001n V_low
+ 591.600000n V_low
+ 591.600001n V_low
+ 591.700000n V_low
+ 591.700001n V_low
+ 591.800000n V_low
+ 591.800001n V_low
+ 591.900000n V_low
+ 591.900001n V_low
+ 592.000000n V_low
+ 592.000001n V_hig
+ 592.100000n V_hig
+ 592.100001n V_hig
+ 592.200000n V_hig
+ 592.200001n V_hig
+ 592.300000n V_hig
+ 592.300001n V_hig
+ 592.400000n V_hig
+ 592.400001n V_hig
+ 592.500000n V_hig
+ 592.500001n V_hig
+ 592.600000n V_hig
+ 592.600001n V_hig
+ 592.700000n V_hig
+ 592.700001n V_hig
+ 592.800000n V_hig
+ 592.800001n V_hig
+ 592.900000n V_hig
+ 592.900001n V_hig
+ 593.000000n V_hig
+ 593.000001n V_hig
+ 593.100000n V_hig
+ 593.100001n V_hig
+ 593.200000n V_hig
+ 593.200001n V_hig
+ 593.300000n V_hig
+ 593.300001n V_hig
+ 593.400000n V_hig
+ 593.400001n V_hig
+ 593.500000n V_hig
+ 593.500001n V_hig
+ 593.600000n V_hig
+ 593.600001n V_hig
+ 593.700000n V_hig
+ 593.700001n V_hig
+ 593.800000n V_hig
+ 593.800001n V_hig
+ 593.900000n V_hig
+ 593.900001n V_hig
+ 594.000000n V_hig
+ 594.000001n V_hig
+ 594.100000n V_hig
+ 594.100001n V_hig
+ 594.200000n V_hig
+ 594.200001n V_hig
+ 594.300000n V_hig
+ 594.300001n V_hig
+ 594.400000n V_hig
+ 594.400001n V_hig
+ 594.500000n V_hig
+ 594.500001n V_hig
+ 594.600000n V_hig
+ 594.600001n V_hig
+ 594.700000n V_hig
+ 594.700001n V_hig
+ 594.800000n V_hig
+ 594.800001n V_hig
+ 594.900000n V_hig
+ 594.900001n V_hig
+ 595.000000n V_hig
+ 595.000001n V_hig
+ 595.100000n V_hig
+ 595.100001n V_hig
+ 595.200000n V_hig
+ 595.200001n V_hig
+ 595.300000n V_hig
+ 595.300001n V_hig
+ 595.400000n V_hig
+ 595.400001n V_hig
+ 595.500000n V_hig
+ 595.500001n V_hig
+ 595.600000n V_hig
+ 595.600001n V_hig
+ 595.700000n V_hig
+ 595.700001n V_hig
+ 595.800000n V_hig
+ 595.800001n V_hig
+ 595.900000n V_hig
+ 595.900001n V_hig
+ 596.000000n V_hig
+ 596.000001n V_hig
+ 596.100000n V_hig
+ 596.100001n V_hig
+ 596.200000n V_hig
+ 596.200001n V_hig
+ 596.300000n V_hig
+ 596.300001n V_hig
+ 596.400000n V_hig
+ 596.400001n V_hig
+ 596.500000n V_hig
+ 596.500001n V_hig
+ 596.600000n V_hig
+ 596.600001n V_hig
+ 596.700000n V_hig
+ 596.700001n V_hig
+ 596.800000n V_hig
+ 596.800001n V_hig
+ 596.900000n V_hig
+ 596.900001n V_hig
+ 597.000000n V_hig
+ 597.000001n V_hig
+ 597.100000n V_hig
+ 597.100001n V_hig
+ 597.200000n V_hig
+ 597.200001n V_hig
+ 597.300000n V_hig
+ 597.300001n V_hig
+ 597.400000n V_hig
+ 597.400001n V_hig
+ 597.500000n V_hig
+ 597.500001n V_hig
+ 597.600000n V_hig
+ 597.600001n V_hig
+ 597.700000n V_hig
+ 597.700001n V_hig
+ 597.800000n V_hig
+ 597.800001n V_hig
+ 597.900000n V_hig
+ 597.900001n V_hig
+ 598.000000n V_hig
+ 598.000001n V_hig
+ 598.100000n V_hig
+ 598.100001n V_hig
+ 598.200000n V_hig
+ 598.200001n V_hig
+ 598.300000n V_hig
+ 598.300001n V_hig
+ 598.400000n V_hig
+ 598.400001n V_hig
+ 598.500000n V_hig
+ 598.500001n V_hig
+ 598.600000n V_hig
+ 598.600001n V_hig
+ 598.700000n V_hig
+ 598.700001n V_hig
+ 598.800000n V_hig
+ 598.800001n V_hig
+ 598.900000n V_hig
+ 598.900001n V_hig
+ 599.000000n V_hig
+ 599.000001n V_low
+ 599.100000n V_low
+ 599.100001n V_low
+ 599.200000n V_low
+ 599.200001n V_low
+ 599.300000n V_low
+ 599.300001n V_low
+ 599.400000n V_low
+ 599.400001n V_low
+ 599.500000n V_low
+ 599.500001n V_low
+ 599.600000n V_low
+ 599.600001n V_low
+ 599.700000n V_low
+ 599.700001n V_low
+ 599.800000n V_low
+ 599.800001n V_low
+ 599.900000n V_low
+ 599.900001n V_low
+ 600.000000n V_low
+ 600.000001n V_hig
+ 600.100000n V_hig
+ 600.100001n V_hig
+ 600.200000n V_hig
+ 600.200001n V_hig
+ 600.300000n V_hig
+ 600.300001n V_hig
+ 600.400000n V_hig
+ 600.400001n V_hig
+ 600.500000n V_hig
+ 600.500001n V_hig
+ 600.600000n V_hig
+ 600.600001n V_hig
+ 600.700000n V_hig
+ 600.700001n V_hig
+ 600.800000n V_hig
+ 600.800001n V_hig
+ 600.900000n V_hig
+ 600.900001n V_hig
+ 601.000000n V_hig
+ 601.000001n V_hig
+ 601.100000n V_hig
+ 601.100001n V_hig
+ 601.200000n V_hig
+ 601.200001n V_hig
+ 601.300000n V_hig
+ 601.300001n V_hig
+ 601.400000n V_hig
+ 601.400001n V_hig
+ 601.500000n V_hig
+ 601.500001n V_hig
+ 601.600000n V_hig
+ 601.600001n V_hig
+ 601.700000n V_hig
+ 601.700001n V_hig
+ 601.800000n V_hig
+ 601.800001n V_hig
+ 601.900000n V_hig
+ 601.900001n V_hig
+ 602.000000n V_hig
+ 602.000001n V_low
+ 602.100000n V_low
+ 602.100001n V_low
+ 602.200000n V_low
+ 602.200001n V_low
+ 602.300000n V_low
+ 602.300001n V_low
+ 602.400000n V_low
+ 602.400001n V_low
+ 602.500000n V_low
+ 602.500001n V_low
+ 602.600000n V_low
+ 602.600001n V_low
+ 602.700000n V_low
+ 602.700001n V_low
+ 602.800000n V_low
+ 602.800001n V_low
+ 602.900000n V_low
+ 602.900001n V_low
+ 603.000000n V_low
+ 603.000001n V_hig
+ 603.100000n V_hig
+ 603.100001n V_hig
+ 603.200000n V_hig
+ 603.200001n V_hig
+ 603.300000n V_hig
+ 603.300001n V_hig
+ 603.400000n V_hig
+ 603.400001n V_hig
+ 603.500000n V_hig
+ 603.500001n V_hig
+ 603.600000n V_hig
+ 603.600001n V_hig
+ 603.700000n V_hig
+ 603.700001n V_hig
+ 603.800000n V_hig
+ 603.800001n V_hig
+ 603.900000n V_hig
+ 603.900001n V_hig
+ 604.000000n V_hig
+ 604.000001n V_hig
+ 604.100000n V_hig
+ 604.100001n V_hig
+ 604.200000n V_hig
+ 604.200001n V_hig
+ 604.300000n V_hig
+ 604.300001n V_hig
+ 604.400000n V_hig
+ 604.400001n V_hig
+ 604.500000n V_hig
+ 604.500001n V_hig
+ 604.600000n V_hig
+ 604.600001n V_hig
+ 604.700000n V_hig
+ 604.700001n V_hig
+ 604.800000n V_hig
+ 604.800001n V_hig
+ 604.900000n V_hig
+ 604.900001n V_hig
+ 605.000000n V_hig
+ 605.000001n V_low
+ 605.100000n V_low
+ 605.100001n V_low
+ 605.200000n V_low
+ 605.200001n V_low
+ 605.300000n V_low
+ 605.300001n V_low
+ 605.400000n V_low
+ 605.400001n V_low
+ 605.500000n V_low
+ 605.500001n V_low
+ 605.600000n V_low
+ 605.600001n V_low
+ 605.700000n V_low
+ 605.700001n V_low
+ 605.800000n V_low
+ 605.800001n V_low
+ 605.900000n V_low
+ 605.900001n V_low
+ 606.000000n V_low
+ 606.000001n V_low
+ 606.100000n V_low
+ 606.100001n V_low
+ 606.200000n V_low
+ 606.200001n V_low
+ 606.300000n V_low
+ 606.300001n V_low
+ 606.400000n V_low
+ 606.400001n V_low
+ 606.500000n V_low
+ 606.500001n V_low
+ 606.600000n V_low
+ 606.600001n V_low
+ 606.700000n V_low
+ 606.700001n V_low
+ 606.800000n V_low
+ 606.800001n V_low
+ 606.900000n V_low
+ 606.900001n V_low
+ 607.000000n V_low
+ 607.000001n V_hig
+ 607.100000n V_hig
+ 607.100001n V_hig
+ 607.200000n V_hig
+ 607.200001n V_hig
+ 607.300000n V_hig
+ 607.300001n V_hig
+ 607.400000n V_hig
+ 607.400001n V_hig
+ 607.500000n V_hig
+ 607.500001n V_hig
+ 607.600000n V_hig
+ 607.600001n V_hig
+ 607.700000n V_hig
+ 607.700001n V_hig
+ 607.800000n V_hig
+ 607.800001n V_hig
+ 607.900000n V_hig
+ 607.900001n V_hig
+ 608.000000n V_hig
+ 608.000001n V_low
+ 608.100000n V_low
+ 608.100001n V_low
+ 608.200000n V_low
+ 608.200001n V_low
+ 608.300000n V_low
+ 608.300001n V_low
+ 608.400000n V_low
+ 608.400001n V_low
+ 608.500000n V_low
+ 608.500001n V_low
+ 608.600000n V_low
+ 608.600001n V_low
+ 608.700000n V_low
+ 608.700001n V_low
+ 608.800000n V_low
+ 608.800001n V_low
+ 608.900000n V_low
+ 608.900001n V_low
+ 609.000000n V_low
+ 609.000001n V_hig
+ 609.100000n V_hig
+ 609.100001n V_hig
+ 609.200000n V_hig
+ 609.200001n V_hig
+ 609.300000n V_hig
+ 609.300001n V_hig
+ 609.400000n V_hig
+ 609.400001n V_hig
+ 609.500000n V_hig
+ 609.500001n V_hig
+ 609.600000n V_hig
+ 609.600001n V_hig
+ 609.700000n V_hig
+ 609.700001n V_hig
+ 609.800000n V_hig
+ 609.800001n V_hig
+ 609.900000n V_hig
+ 609.900001n V_hig
+ 610.000000n V_hig
+ 610.000001n V_hig
+ 610.100000n V_hig
+ 610.100001n V_hig
+ 610.200000n V_hig
+ 610.200001n V_hig
+ 610.300000n V_hig
+ 610.300001n V_hig
+ 610.400000n V_hig
+ 610.400001n V_hig
+ 610.500000n V_hig
+ 610.500001n V_hig
+ 610.600000n V_hig
+ 610.600001n V_hig
+ 610.700000n V_hig
+ 610.700001n V_hig
+ 610.800000n V_hig
+ 610.800001n V_hig
+ 610.900000n V_hig
+ 610.900001n V_hig
+ 611.000000n V_hig
+ 611.000001n V_low
+ 611.100000n V_low
+ 611.100001n V_low
+ 611.200000n V_low
+ 611.200001n V_low
+ 611.300000n V_low
+ 611.300001n V_low
+ 611.400000n V_low
+ 611.400001n V_low
+ 611.500000n V_low
+ 611.500001n V_low
+ 611.600000n V_low
+ 611.600001n V_low
+ 611.700000n V_low
+ 611.700001n V_low
+ 611.800000n V_low
+ 611.800001n V_low
+ 611.900000n V_low
+ 611.900001n V_low
+ 612.000000n V_low
+ 612.000001n V_low
+ 612.100000n V_low
+ 612.100001n V_low
+ 612.200000n V_low
+ 612.200001n V_low
+ 612.300000n V_low
+ 612.300001n V_low
+ 612.400000n V_low
+ 612.400001n V_low
+ 612.500000n V_low
+ 612.500001n V_low
+ 612.600000n V_low
+ 612.600001n V_low
+ 612.700000n V_low
+ 612.700001n V_low
+ 612.800000n V_low
+ 612.800001n V_low
+ 612.900000n V_low
+ 612.900001n V_low
+ 613.000000n V_low
+ 613.000001n V_hig
+ 613.100000n V_hig
+ 613.100001n V_hig
+ 613.200000n V_hig
+ 613.200001n V_hig
+ 613.300000n V_hig
+ 613.300001n V_hig
+ 613.400000n V_hig
+ 613.400001n V_hig
+ 613.500000n V_hig
+ 613.500001n V_hig
+ 613.600000n V_hig
+ 613.600001n V_hig
+ 613.700000n V_hig
+ 613.700001n V_hig
+ 613.800000n V_hig
+ 613.800001n V_hig
+ 613.900000n V_hig
+ 613.900001n V_hig
+ 614.000000n V_hig
+ 614.000001n V_low
+ 614.100000n V_low
+ 614.100001n V_low
+ 614.200000n V_low
+ 614.200001n V_low
+ 614.300000n V_low
+ 614.300001n V_low
+ 614.400000n V_low
+ 614.400001n V_low
+ 614.500000n V_low
+ 614.500001n V_low
+ 614.600000n V_low
+ 614.600001n V_low
+ 614.700000n V_low
+ 614.700001n V_low
+ 614.800000n V_low
+ 614.800001n V_low
+ 614.900000n V_low
+ 614.900001n V_low
+ 615.000000n V_low
+ 615.000001n V_hig
+ 615.100000n V_hig
+ 615.100001n V_hig
+ 615.200000n V_hig
+ 615.200001n V_hig
+ 615.300000n V_hig
+ 615.300001n V_hig
+ 615.400000n V_hig
+ 615.400001n V_hig
+ 615.500000n V_hig
+ 615.500001n V_hig
+ 615.600000n V_hig
+ 615.600001n V_hig
+ 615.700000n V_hig
+ 615.700001n V_hig
+ 615.800000n V_hig
+ 615.800001n V_hig
+ 615.900000n V_hig
+ 615.900001n V_hig
+ 616.000000n V_hig
+ 616.000001n V_low
+ 616.100000n V_low
+ 616.100001n V_low
+ 616.200000n V_low
+ 616.200001n V_low
+ 616.300000n V_low
+ 616.300001n V_low
+ 616.400000n V_low
+ 616.400001n V_low
+ 616.500000n V_low
+ 616.500001n V_low
+ 616.600000n V_low
+ 616.600001n V_low
+ 616.700000n V_low
+ 616.700001n V_low
+ 616.800000n V_low
+ 616.800001n V_low
+ 616.900000n V_low
+ 616.900001n V_low
+ 617.000000n V_low
+ 617.000001n V_low
+ 617.100000n V_low
+ 617.100001n V_low
+ 617.200000n V_low
+ 617.200001n V_low
+ 617.300000n V_low
+ 617.300001n V_low
+ 617.400000n V_low
+ 617.400001n V_low
+ 617.500000n V_low
+ 617.500001n V_low
+ 617.600000n V_low
+ 617.600001n V_low
+ 617.700000n V_low
+ 617.700001n V_low
+ 617.800000n V_low
+ 617.800001n V_low
+ 617.900000n V_low
+ 617.900001n V_low
+ 618.000000n V_low
+ 618.000001n V_low
+ 618.100000n V_low
+ 618.100001n V_low
+ 618.200000n V_low
+ 618.200001n V_low
+ 618.300000n V_low
+ 618.300001n V_low
+ 618.400000n V_low
+ 618.400001n V_low
+ 618.500000n V_low
+ 618.500001n V_low
+ 618.600000n V_low
+ 618.600001n V_low
+ 618.700000n V_low
+ 618.700001n V_low
+ 618.800000n V_low
+ 618.800001n V_low
+ 618.900000n V_low
+ 618.900001n V_low
+ 619.000000n V_low
+ 619.000001n V_hig
+ 619.100000n V_hig
+ 619.100001n V_hig
+ 619.200000n V_hig
+ 619.200001n V_hig
+ 619.300000n V_hig
+ 619.300001n V_hig
+ 619.400000n V_hig
+ 619.400001n V_hig
+ 619.500000n V_hig
+ 619.500001n V_hig
+ 619.600000n V_hig
+ 619.600001n V_hig
+ 619.700000n V_hig
+ 619.700001n V_hig
+ 619.800000n V_hig
+ 619.800001n V_hig
+ 619.900000n V_hig
+ 619.900001n V_hig
+ 620.000000n V_hig
+ 620.000001n V_low
+ 620.100000n V_low
+ 620.100001n V_low
+ 620.200000n V_low
+ 620.200001n V_low
+ 620.300000n V_low
+ 620.300001n V_low
+ 620.400000n V_low
+ 620.400001n V_low
+ 620.500000n V_low
+ 620.500001n V_low
+ 620.600000n V_low
+ 620.600001n V_low
+ 620.700000n V_low
+ 620.700001n V_low
+ 620.800000n V_low
+ 620.800001n V_low
+ 620.900000n V_low
+ 620.900001n V_low
+ 621.000000n V_low
+ 621.000001n V_hig
+ 621.100000n V_hig
+ 621.100001n V_hig
+ 621.200000n V_hig
+ 621.200001n V_hig
+ 621.300000n V_hig
+ 621.300001n V_hig
+ 621.400000n V_hig
+ 621.400001n V_hig
+ 621.500000n V_hig
+ 621.500001n V_hig
+ 621.600000n V_hig
+ 621.600001n V_hig
+ 621.700000n V_hig
+ 621.700001n V_hig
+ 621.800000n V_hig
+ 621.800001n V_hig
+ 621.900000n V_hig
+ 621.900001n V_hig
+ 622.000000n V_hig
+ 622.000001n V_low
+ 622.100000n V_low
+ 622.100001n V_low
+ 622.200000n V_low
+ 622.200001n V_low
+ 622.300000n V_low
+ 622.300001n V_low
+ 622.400000n V_low
+ 622.400001n V_low
+ 622.500000n V_low
+ 622.500001n V_low
+ 622.600000n V_low
+ 622.600001n V_low
+ 622.700000n V_low
+ 622.700001n V_low
+ 622.800000n V_low
+ 622.800001n V_low
+ 622.900000n V_low
+ 622.900001n V_low
+ 623.000000n V_low
+ 623.000001n V_hig
+ 623.100000n V_hig
+ 623.100001n V_hig
+ 623.200000n V_hig
+ 623.200001n V_hig
+ 623.300000n V_hig
+ 623.300001n V_hig
+ 623.400000n V_hig
+ 623.400001n V_hig
+ 623.500000n V_hig
+ 623.500001n V_hig
+ 623.600000n V_hig
+ 623.600001n V_hig
+ 623.700000n V_hig
+ 623.700001n V_hig
+ 623.800000n V_hig
+ 623.800001n V_hig
+ 623.900000n V_hig
+ 623.900001n V_hig
+ 624.000000n V_hig
+ 624.000001n V_low
+ 624.100000n V_low
+ 624.100001n V_low
+ 624.200000n V_low
+ 624.200001n V_low
+ 624.300000n V_low
+ 624.300001n V_low
+ 624.400000n V_low
+ 624.400001n V_low
+ 624.500000n V_low
+ 624.500001n V_low
+ 624.600000n V_low
+ 624.600001n V_low
+ 624.700000n V_low
+ 624.700001n V_low
+ 624.800000n V_low
+ 624.800001n V_low
+ 624.900000n V_low
+ 624.900001n V_low
+ 625.000000n V_low
+ 625.000001n V_low
+ 625.100000n V_low
+ 625.100001n V_low
+ 625.200000n V_low
+ 625.200001n V_low
+ 625.300000n V_low
+ 625.300001n V_low
+ 625.400000n V_low
+ 625.400001n V_low
+ 625.500000n V_low
+ 625.500001n V_low
+ 625.600000n V_low
+ 625.600001n V_low
+ 625.700000n V_low
+ 625.700001n V_low
+ 625.800000n V_low
+ 625.800001n V_low
+ 625.900000n V_low
+ 625.900001n V_low
+ 626.000000n V_low
+ 626.000001n V_low
+ 626.100000n V_low
+ 626.100001n V_low
+ 626.200000n V_low
+ 626.200001n V_low
+ 626.300000n V_low
+ 626.300001n V_low
+ 626.400000n V_low
+ 626.400001n V_low
+ 626.500000n V_low
+ 626.500001n V_low
+ 626.600000n V_low
+ 626.600001n V_low
+ 626.700000n V_low
+ 626.700001n V_low
+ 626.800000n V_low
+ 626.800001n V_low
+ 626.900000n V_low
+ 626.900001n V_low
+ 627.000000n V_low
+ 627.000001n V_low
+ 627.100000n V_low
+ 627.100001n V_low
+ 627.200000n V_low
+ 627.200001n V_low
+ 627.300000n V_low
+ 627.300001n V_low
+ 627.400000n V_low
+ 627.400001n V_low
+ 627.500000n V_low
+ 627.500001n V_low
+ 627.600000n V_low
+ 627.600001n V_low
+ 627.700000n V_low
+ 627.700001n V_low
+ 627.800000n V_low
+ 627.800001n V_low
+ 627.900000n V_low
+ 627.900001n V_low
+ 628.000000n V_low
+ 628.000001n V_low
+ 628.100000n V_low
+ 628.100001n V_low
+ 628.200000n V_low
+ 628.200001n V_low
+ 628.300000n V_low
+ 628.300001n V_low
+ 628.400000n V_low
+ 628.400001n V_low
+ 628.500000n V_low
+ 628.500001n V_low
+ 628.600000n V_low
+ 628.600001n V_low
+ 628.700000n V_low
+ 628.700001n V_low
+ 628.800000n V_low
+ 628.800001n V_low
+ 628.900000n V_low
+ 628.900001n V_low
+ 629.000000n V_low
+ 629.000001n V_low
+ 629.100000n V_low
+ 629.100001n V_low
+ 629.200000n V_low
+ 629.200001n V_low
+ 629.300000n V_low
+ 629.300001n V_low
+ 629.400000n V_low
+ 629.400001n V_low
+ 629.500000n V_low
+ 629.500001n V_low
+ 629.600000n V_low
+ 629.600001n V_low
+ 629.700000n V_low
+ 629.700001n V_low
+ 629.800000n V_low
+ 629.800001n V_low
+ 629.900000n V_low
+ 629.900001n V_low
+ 630.000000n V_low
+ 630.000001n V_low
+ 630.100000n V_low
+ 630.100001n V_low
+ 630.200000n V_low
+ 630.200001n V_low
+ 630.300000n V_low
+ 630.300001n V_low
+ 630.400000n V_low
+ 630.400001n V_low
+ 630.500000n V_low
+ 630.500001n V_low
+ 630.600000n V_low
+ 630.600001n V_low
+ 630.700000n V_low
+ 630.700001n V_low
+ 630.800000n V_low
+ 630.800001n V_low
+ 630.900000n V_low
+ 630.900001n V_low
+ 631.000000n V_low
+ 631.000001n V_hig
+ 631.100000n V_hig
+ 631.100001n V_hig
+ 631.200000n V_hig
+ 631.200001n V_hig
+ 631.300000n V_hig
+ 631.300001n V_hig
+ 631.400000n V_hig
+ 631.400001n V_hig
+ 631.500000n V_hig
+ 631.500001n V_hig
+ 631.600000n V_hig
+ 631.600001n V_hig
+ 631.700000n V_hig
+ 631.700001n V_hig
+ 631.800000n V_hig
+ 631.800001n V_hig
+ 631.900000n V_hig
+ 631.900001n V_hig
+ 632.000000n V_hig
+ 632.000001n V_low
+ 632.100000n V_low
+ 632.100001n V_low
+ 632.200000n V_low
+ 632.200001n V_low
+ 632.300000n V_low
+ 632.300001n V_low
+ 632.400000n V_low
+ 632.400001n V_low
+ 632.500000n V_low
+ 632.500001n V_low
+ 632.600000n V_low
+ 632.600001n V_low
+ 632.700000n V_low
+ 632.700001n V_low
+ 632.800000n V_low
+ 632.800001n V_low
+ 632.900000n V_low
+ 632.900001n V_low
+ 633.000000n V_low
+ 633.000001n V_low
+ 633.100000n V_low
+ 633.100001n V_low
+ 633.200000n V_low
+ 633.200001n V_low
+ 633.300000n V_low
+ 633.300001n V_low
+ 633.400000n V_low
+ 633.400001n V_low
+ 633.500000n V_low
+ 633.500001n V_low
+ 633.600000n V_low
+ 633.600001n V_low
+ 633.700000n V_low
+ 633.700001n V_low
+ 633.800000n V_low
+ 633.800001n V_low
+ 633.900000n V_low
+ 633.900001n V_low
+ 634.000000n V_low
+ 634.000001n V_low
+ 634.100000n V_low
+ 634.100001n V_low
+ 634.200000n V_low
+ 634.200001n V_low
+ 634.300000n V_low
+ 634.300001n V_low
+ 634.400000n V_low
+ 634.400001n V_low
+ 634.500000n V_low
+ 634.500001n V_low
+ 634.600000n V_low
+ 634.600001n V_low
+ 634.700000n V_low
+ 634.700001n V_low
+ 634.800000n V_low
+ 634.800001n V_low
+ 634.900000n V_low
+ 634.900001n V_low
+ 635.000000n V_low
+ 635.000001n V_hig
+ 635.100000n V_hig
+ 635.100001n V_hig
+ 635.200000n V_hig
+ 635.200001n V_hig
+ 635.300000n V_hig
+ 635.300001n V_hig
+ 635.400000n V_hig
+ 635.400001n V_hig
+ 635.500000n V_hig
+ 635.500001n V_hig
+ 635.600000n V_hig
+ 635.600001n V_hig
+ 635.700000n V_hig
+ 635.700001n V_hig
+ 635.800000n V_hig
+ 635.800001n V_hig
+ 635.900000n V_hig
+ 635.900001n V_hig
+ 636.000000n V_hig
+ 636.000001n V_low
+ 636.100000n V_low
+ 636.100001n V_low
+ 636.200000n V_low
+ 636.200001n V_low
+ 636.300000n V_low
+ 636.300001n V_low
+ 636.400000n V_low
+ 636.400001n V_low
+ 636.500000n V_low
+ 636.500001n V_low
+ 636.600000n V_low
+ 636.600001n V_low
+ 636.700000n V_low
+ 636.700001n V_low
+ 636.800000n V_low
+ 636.800001n V_low
+ 636.900000n V_low
+ 636.900001n V_low
+ 637.000000n V_low
+ 637.000001n V_low
+ 637.100000n V_low
+ 637.100001n V_low
+ 637.200000n V_low
+ 637.200001n V_low
+ 637.300000n V_low
+ 637.300001n V_low
+ 637.400000n V_low
+ 637.400001n V_low
+ 637.500000n V_low
+ 637.500001n V_low
+ 637.600000n V_low
+ 637.600001n V_low
+ 637.700000n V_low
+ 637.700001n V_low
+ 637.800000n V_low
+ 637.800001n V_low
+ 637.900000n V_low
+ 637.900001n V_low
+ 638.000000n V_low
+ 638.000001n V_hig
+ 638.100000n V_hig
+ 638.100001n V_hig
+ 638.200000n V_hig
+ 638.200001n V_hig
+ 638.300000n V_hig
+ 638.300001n V_hig
+ 638.400000n V_hig
+ 638.400001n V_hig
+ 638.500000n V_hig
+ 638.500001n V_hig
+ 638.600000n V_hig
+ 638.600001n V_hig
+ 638.700000n V_hig
+ 638.700001n V_hig
+ 638.800000n V_hig
+ 638.800001n V_hig
+ 638.900000n V_hig
+ 638.900001n V_hig
+ 639.000000n V_hig
+ 639.000001n V_low
+ 639.100000n V_low
+ 639.100001n V_low
+ 639.200000n V_low
+ 639.200001n V_low
+ 639.300000n V_low
+ 639.300001n V_low
+ 639.400000n V_low
+ 639.400001n V_low
+ 639.500000n V_low
+ 639.500001n V_low
+ 639.600000n V_low
+ 639.600001n V_low
+ 639.700000n V_low
+ 639.700001n V_low
+ 639.800000n V_low
+ 639.800001n V_low
+ 639.900000n V_low
+ 639.900001n V_low
+ 640.000000n V_low
+ 640.000001n V_low
+ 640.100000n V_low
+ 640.100001n V_low
+ 640.200000n V_low
+ 640.200001n V_low
+ 640.300000n V_low
+ 640.300001n V_low
+ 640.400000n V_low
+ 640.400001n V_low
+ 640.500000n V_low
+ 640.500001n V_low
+ 640.600000n V_low
+ 640.600001n V_low
+ 640.700000n V_low
+ 640.700001n V_low
+ 640.800000n V_low
+ 640.800001n V_low
+ 640.900000n V_low
+ 640.900001n V_low
+ 641.000000n V_low
+ 641.000001n V_low
+ 641.100000n V_low
+ 641.100001n V_low
+ 641.200000n V_low
+ 641.200001n V_low
+ 641.300000n V_low
+ 641.300001n V_low
+ 641.400000n V_low
+ 641.400001n V_low
+ 641.500000n V_low
+ 641.500001n V_low
+ 641.600000n V_low
+ 641.600001n V_low
+ 641.700000n V_low
+ 641.700001n V_low
+ 641.800000n V_low
+ 641.800001n V_low
+ 641.900000n V_low
+ 641.900001n V_low
+ 642.000000n V_low
+ 642.000001n V_low
+ 642.100000n V_low
+ 642.100001n V_low
+ 642.200000n V_low
+ 642.200001n V_low
+ 642.300000n V_low
+ 642.300001n V_low
+ 642.400000n V_low
+ 642.400001n V_low
+ 642.500000n V_low
+ 642.500001n V_low
+ 642.600000n V_low
+ 642.600001n V_low
+ 642.700000n V_low
+ 642.700001n V_low
+ 642.800000n V_low
+ 642.800001n V_low
+ 642.900000n V_low
+ 642.900001n V_low
+ 643.000000n V_low
+ 643.000001n V_hig
+ 643.100000n V_hig
+ 643.100001n V_hig
+ 643.200000n V_hig
+ 643.200001n V_hig
+ 643.300000n V_hig
+ 643.300001n V_hig
+ 643.400000n V_hig
+ 643.400001n V_hig
+ 643.500000n V_hig
+ 643.500001n V_hig
+ 643.600000n V_hig
+ 643.600001n V_hig
+ 643.700000n V_hig
+ 643.700001n V_hig
+ 643.800000n V_hig
+ 643.800001n V_hig
+ 643.900000n V_hig
+ 643.900001n V_hig
+ 644.000000n V_hig
+ 644.000001n V_low
+ 644.100000n V_low
+ 644.100001n V_low
+ 644.200000n V_low
+ 644.200001n V_low
+ 644.300000n V_low
+ 644.300001n V_low
+ 644.400000n V_low
+ 644.400001n V_low
+ 644.500000n V_low
+ 644.500001n V_low
+ 644.600000n V_low
+ 644.600001n V_low
+ 644.700000n V_low
+ 644.700001n V_low
+ 644.800000n V_low
+ 644.800001n V_low
+ 644.900000n V_low
+ 644.900001n V_low
+ 645.000000n V_low
+ 645.000001n V_low
+ 645.100000n V_low
+ 645.100001n V_low
+ 645.200000n V_low
+ 645.200001n V_low
+ 645.300000n V_low
+ 645.300001n V_low
+ 645.400000n V_low
+ 645.400001n V_low
+ 645.500000n V_low
+ 645.500001n V_low
+ 645.600000n V_low
+ 645.600001n V_low
+ 645.700000n V_low
+ 645.700001n V_low
+ 645.800000n V_low
+ 645.800001n V_low
+ 645.900000n V_low
+ 645.900001n V_low
+ 646.000000n V_low
+ 646.000001n V_hig
+ 646.100000n V_hig
+ 646.100001n V_hig
+ 646.200000n V_hig
+ 646.200001n V_hig
+ 646.300000n V_hig
+ 646.300001n V_hig
+ 646.400000n V_hig
+ 646.400001n V_hig
+ 646.500000n V_hig
+ 646.500001n V_hig
+ 646.600000n V_hig
+ 646.600001n V_hig
+ 646.700000n V_hig
+ 646.700001n V_hig
+ 646.800000n V_hig
+ 646.800001n V_hig
+ 646.900000n V_hig
+ 646.900001n V_hig
+ 647.000000n V_hig
+ 647.000001n V_hig
+ 647.100000n V_hig
+ 647.100001n V_hig
+ 647.200000n V_hig
+ 647.200001n V_hig
+ 647.300000n V_hig
+ 647.300001n V_hig
+ 647.400000n V_hig
+ 647.400001n V_hig
+ 647.500000n V_hig
+ 647.500001n V_hig
+ 647.600000n V_hig
+ 647.600001n V_hig
+ 647.700000n V_hig
+ 647.700001n V_hig
+ 647.800000n V_hig
+ 647.800001n V_hig
+ 647.900000n V_hig
+ 647.900001n V_hig
+ 648.000000n V_hig
+ 648.000001n V_low
+ 648.100000n V_low
+ 648.100001n V_low
+ 648.200000n V_low
+ 648.200001n V_low
+ 648.300000n V_low
+ 648.300001n V_low
+ 648.400000n V_low
+ 648.400001n V_low
+ 648.500000n V_low
+ 648.500001n V_low
+ 648.600000n V_low
+ 648.600001n V_low
+ 648.700000n V_low
+ 648.700001n V_low
+ 648.800000n V_low
+ 648.800001n V_low
+ 648.900000n V_low
+ 648.900001n V_low
+ 649.000000n V_low
+ 649.000001n V_low
+ 649.100000n V_low
+ 649.100001n V_low
+ 649.200000n V_low
+ 649.200001n V_low
+ 649.300000n V_low
+ 649.300001n V_low
+ 649.400000n V_low
+ 649.400001n V_low
+ 649.500000n V_low
+ 649.500001n V_low
+ 649.600000n V_low
+ 649.600001n V_low
+ 649.700000n V_low
+ 649.700001n V_low
+ 649.800000n V_low
+ 649.800001n V_low
+ 649.900000n V_low
+ 649.900001n V_low
+ 650.000000n V_low
+ 650.000001n V_hig
+ 650.100000n V_hig
+ 650.100001n V_hig
+ 650.200000n V_hig
+ 650.200001n V_hig
+ 650.300000n V_hig
+ 650.300001n V_hig
+ 650.400000n V_hig
+ 650.400001n V_hig
+ 650.500000n V_hig
+ 650.500001n V_hig
+ 650.600000n V_hig
+ 650.600001n V_hig
+ 650.700000n V_hig
+ 650.700001n V_hig
+ 650.800000n V_hig
+ 650.800001n V_hig
+ 650.900000n V_hig
+ 650.900001n V_hig
+ 651.000000n V_hig
+ 651.000001n V_hig
+ 651.100000n V_hig
+ 651.100001n V_hig
+ 651.200000n V_hig
+ 651.200001n V_hig
+ 651.300000n V_hig
+ 651.300001n V_hig
+ 651.400000n V_hig
+ 651.400001n V_hig
+ 651.500000n V_hig
+ 651.500001n V_hig
+ 651.600000n V_hig
+ 651.600001n V_hig
+ 651.700000n V_hig
+ 651.700001n V_hig
+ 651.800000n V_hig
+ 651.800001n V_hig
+ 651.900000n V_hig
+ 651.900001n V_hig
+ 652.000000n V_hig
+ 652.000001n V_low
+ 652.100000n V_low
+ 652.100001n V_low
+ 652.200000n V_low
+ 652.200001n V_low
+ 652.300000n V_low
+ 652.300001n V_low
+ 652.400000n V_low
+ 652.400001n V_low
+ 652.500000n V_low
+ 652.500001n V_low
+ 652.600000n V_low
+ 652.600001n V_low
+ 652.700000n V_low
+ 652.700001n V_low
+ 652.800000n V_low
+ 652.800001n V_low
+ 652.900000n V_low
+ 652.900001n V_low
+ 653.000000n V_low
+ 653.000001n V_low
+ 653.100000n V_low
+ 653.100001n V_low
+ 653.200000n V_low
+ 653.200001n V_low
+ 653.300000n V_low
+ 653.300001n V_low
+ 653.400000n V_low
+ 653.400001n V_low
+ 653.500000n V_low
+ 653.500001n V_low
+ 653.600000n V_low
+ 653.600001n V_low
+ 653.700000n V_low
+ 653.700001n V_low
+ 653.800000n V_low
+ 653.800001n V_low
+ 653.900000n V_low
+ 653.900001n V_low
+ 654.000000n V_low
+ 654.000001n V_hig
+ 654.100000n V_hig
+ 654.100001n V_hig
+ 654.200000n V_hig
+ 654.200001n V_hig
+ 654.300000n V_hig
+ 654.300001n V_hig
+ 654.400000n V_hig
+ 654.400001n V_hig
+ 654.500000n V_hig
+ 654.500001n V_hig
+ 654.600000n V_hig
+ 654.600001n V_hig
+ 654.700000n V_hig
+ 654.700001n V_hig
+ 654.800000n V_hig
+ 654.800001n V_hig
+ 654.900000n V_hig
+ 654.900001n V_hig
+ 655.000000n V_hig
+ 655.000001n V_hig
+ 655.100000n V_hig
+ 655.100001n V_hig
+ 655.200000n V_hig
+ 655.200001n V_hig
+ 655.300000n V_hig
+ 655.300001n V_hig
+ 655.400000n V_hig
+ 655.400001n V_hig
+ 655.500000n V_hig
+ 655.500001n V_hig
+ 655.600000n V_hig
+ 655.600001n V_hig
+ 655.700000n V_hig
+ 655.700001n V_hig
+ 655.800000n V_hig
+ 655.800001n V_hig
+ 655.900000n V_hig
+ 655.900001n V_hig
+ 656.000000n V_hig
+ 656.000001n V_hig
+ 656.100000n V_hig
+ 656.100001n V_hig
+ 656.200000n V_hig
+ 656.200001n V_hig
+ 656.300000n V_hig
+ 656.300001n V_hig
+ 656.400000n V_hig
+ 656.400001n V_hig
+ 656.500000n V_hig
+ 656.500001n V_hig
+ 656.600000n V_hig
+ 656.600001n V_hig
+ 656.700000n V_hig
+ 656.700001n V_hig
+ 656.800000n V_hig
+ 656.800001n V_hig
+ 656.900000n V_hig
+ 656.900001n V_hig
+ 657.000000n V_hig
+ 657.000001n V_hig
+ 657.100000n V_hig
+ 657.100001n V_hig
+ 657.200000n V_hig
+ 657.200001n V_hig
+ 657.300000n V_hig
+ 657.300001n V_hig
+ 657.400000n V_hig
+ 657.400001n V_hig
+ 657.500000n V_hig
+ 657.500001n V_hig
+ 657.600000n V_hig
+ 657.600001n V_hig
+ 657.700000n V_hig
+ 657.700001n V_hig
+ 657.800000n V_hig
+ 657.800001n V_hig
+ 657.900000n V_hig
+ 657.900001n V_hig
+ 658.000000n V_hig
+ 658.000001n V_hig
+ 658.100000n V_hig
+ 658.100001n V_hig
+ 658.200000n V_hig
+ 658.200001n V_hig
+ 658.300000n V_hig
+ 658.300001n V_hig
+ 658.400000n V_hig
+ 658.400001n V_hig
+ 658.500000n V_hig
+ 658.500001n V_hig
+ 658.600000n V_hig
+ 658.600001n V_hig
+ 658.700000n V_hig
+ 658.700001n V_hig
+ 658.800000n V_hig
+ 658.800001n V_hig
+ 658.900000n V_hig
+ 658.900001n V_hig
+ 659.000000n V_hig
+ 659.000001n V_hig
+ 659.100000n V_hig
+ 659.100001n V_hig
+ 659.200000n V_hig
+ 659.200001n V_hig
+ 659.300000n V_hig
+ 659.300001n V_hig
+ 659.400000n V_hig
+ 659.400001n V_hig
+ 659.500000n V_hig
+ 659.500001n V_hig
+ 659.600000n V_hig
+ 659.600001n V_hig
+ 659.700000n V_hig
+ 659.700001n V_hig
+ 659.800000n V_hig
+ 659.800001n V_hig
+ 659.900000n V_hig
+ 659.900001n V_hig
+ 660.000000n V_hig
+ 660.000001n V_low
+ 660.100000n V_low
+ 660.100001n V_low
+ 660.200000n V_low
+ 660.200001n V_low
+ 660.300000n V_low
+ 660.300001n V_low
+ 660.400000n V_low
+ 660.400001n V_low
+ 660.500000n V_low
+ 660.500001n V_low
+ 660.600000n V_low
+ 660.600001n V_low
+ 660.700000n V_low
+ 660.700001n V_low
+ 660.800000n V_low
+ 660.800001n V_low
+ 660.900000n V_low
+ 660.900001n V_low
+ 661.000000n V_low
+ 661.000001n V_low
+ 661.100000n V_low
+ 661.100001n V_low
+ 661.200000n V_low
+ 661.200001n V_low
+ 661.300000n V_low
+ 661.300001n V_low
+ 661.400000n V_low
+ 661.400001n V_low
+ 661.500000n V_low
+ 661.500001n V_low
+ 661.600000n V_low
+ 661.600001n V_low
+ 661.700000n V_low
+ 661.700001n V_low
+ 661.800000n V_low
+ 661.800001n V_low
+ 661.900000n V_low
+ 661.900001n V_low
+ 662.000000n V_low
+ 662.000001n V_low
+ 662.100000n V_low
+ 662.100001n V_low
+ 662.200000n V_low
+ 662.200001n V_low
+ 662.300000n V_low
+ 662.300001n V_low
+ 662.400000n V_low
+ 662.400001n V_low
+ 662.500000n V_low
+ 662.500001n V_low
+ 662.600000n V_low
+ 662.600001n V_low
+ 662.700000n V_low
+ 662.700001n V_low
+ 662.800000n V_low
+ 662.800001n V_low
+ 662.900000n V_low
+ 662.900001n V_low
+ 663.000000n V_low
+ 663.000001n V_hig
+ 663.100000n V_hig
+ 663.100001n V_hig
+ 663.200000n V_hig
+ 663.200001n V_hig
+ 663.300000n V_hig
+ 663.300001n V_hig
+ 663.400000n V_hig
+ 663.400001n V_hig
+ 663.500000n V_hig
+ 663.500001n V_hig
+ 663.600000n V_hig
+ 663.600001n V_hig
+ 663.700000n V_hig
+ 663.700001n V_hig
+ 663.800000n V_hig
+ 663.800001n V_hig
+ 663.900000n V_hig
+ 663.900001n V_hig
+ 664.000000n V_hig
+ 664.000001n V_low
+ 664.100000n V_low
+ 664.100001n V_low
+ 664.200000n V_low
+ 664.200001n V_low
+ 664.300000n V_low
+ 664.300001n V_low
+ 664.400000n V_low
+ 664.400001n V_low
+ 664.500000n V_low
+ 664.500001n V_low
+ 664.600000n V_low
+ 664.600001n V_low
+ 664.700000n V_low
+ 664.700001n V_low
+ 664.800000n V_low
+ 664.800001n V_low
+ 664.900000n V_low
+ 664.900001n V_low
+ 665.000000n V_low
+ 665.000001n V_low
+ 665.100000n V_low
+ 665.100001n V_low
+ 665.200000n V_low
+ 665.200001n V_low
+ 665.300000n V_low
+ 665.300001n V_low
+ 665.400000n V_low
+ 665.400001n V_low
+ 665.500000n V_low
+ 665.500001n V_low
+ 665.600000n V_low
+ 665.600001n V_low
+ 665.700000n V_low
+ 665.700001n V_low
+ 665.800000n V_low
+ 665.800001n V_low
+ 665.900000n V_low
+ 665.900001n V_low
+ 666.000000n V_low
+ 666.000001n V_low
+ 666.100000n V_low
+ 666.100001n V_low
+ 666.200000n V_low
+ 666.200001n V_low
+ 666.300000n V_low
+ 666.300001n V_low
+ 666.400000n V_low
+ 666.400001n V_low
+ 666.500000n V_low
+ 666.500001n V_low
+ 666.600000n V_low
+ 666.600001n V_low
+ 666.700000n V_low
+ 666.700001n V_low
+ 666.800000n V_low
+ 666.800001n V_low
+ 666.900000n V_low
+ 666.900001n V_low
+ 667.000000n V_low
+ 667.000001n V_hig
+ 667.100000n V_hig
+ 667.100001n V_hig
+ 667.200000n V_hig
+ 667.200001n V_hig
+ 667.300000n V_hig
+ 667.300001n V_hig
+ 667.400000n V_hig
+ 667.400001n V_hig
+ 667.500000n V_hig
+ 667.500001n V_hig
+ 667.600000n V_hig
+ 667.600001n V_hig
+ 667.700000n V_hig
+ 667.700001n V_hig
+ 667.800000n V_hig
+ 667.800001n V_hig
+ 667.900000n V_hig
+ 667.900001n V_hig
+ 668.000000n V_hig
+ 668.000001n V_hig
+ 668.100000n V_hig
+ 668.100001n V_hig
+ 668.200000n V_hig
+ 668.200001n V_hig
+ 668.300000n V_hig
+ 668.300001n V_hig
+ 668.400000n V_hig
+ 668.400001n V_hig
+ 668.500000n V_hig
+ 668.500001n V_hig
+ 668.600000n V_hig
+ 668.600001n V_hig
+ 668.700000n V_hig
+ 668.700001n V_hig
+ 668.800000n V_hig
+ 668.800001n V_hig
+ 668.900000n V_hig
+ 668.900001n V_hig
+ 669.000000n V_hig
+ 669.000001n V_hig
+ 669.100000n V_hig
+ 669.100001n V_hig
+ 669.200000n V_hig
+ 669.200001n V_hig
+ 669.300000n V_hig
+ 669.300001n V_hig
+ 669.400000n V_hig
+ 669.400001n V_hig
+ 669.500000n V_hig
+ 669.500001n V_hig
+ 669.600000n V_hig
+ 669.600001n V_hig
+ 669.700000n V_hig
+ 669.700001n V_hig
+ 669.800000n V_hig
+ 669.800001n V_hig
+ 669.900000n V_hig
+ 669.900001n V_hig
+ 670.000000n V_hig
+ 670.000001n V_low
+ 670.100000n V_low
+ 670.100001n V_low
+ 670.200000n V_low
+ 670.200001n V_low
+ 670.300000n V_low
+ 670.300001n V_low
+ 670.400000n V_low
+ 670.400001n V_low
+ 670.500000n V_low
+ 670.500001n V_low
+ 670.600000n V_low
+ 670.600001n V_low
+ 670.700000n V_low
+ 670.700001n V_low
+ 670.800000n V_low
+ 670.800001n V_low
+ 670.900000n V_low
+ 670.900001n V_low
+ 671.000000n V_low
+ 671.000001n V_hig
+ 671.100000n V_hig
+ 671.100001n V_hig
+ 671.200000n V_hig
+ 671.200001n V_hig
+ 671.300000n V_hig
+ 671.300001n V_hig
+ 671.400000n V_hig
+ 671.400001n V_hig
+ 671.500000n V_hig
+ 671.500001n V_hig
+ 671.600000n V_hig
+ 671.600001n V_hig
+ 671.700000n V_hig
+ 671.700001n V_hig
+ 671.800000n V_hig
+ 671.800001n V_hig
+ 671.900000n V_hig
+ 671.900001n V_hig
+ 672.000000n V_hig
+ 672.000001n V_hig
+ 672.100000n V_hig
+ 672.100001n V_hig
+ 672.200000n V_hig
+ 672.200001n V_hig
+ 672.300000n V_hig
+ 672.300001n V_hig
+ 672.400000n V_hig
+ 672.400001n V_hig
+ 672.500000n V_hig
+ 672.500001n V_hig
+ 672.600000n V_hig
+ 672.600001n V_hig
+ 672.700000n V_hig
+ 672.700001n V_hig
+ 672.800000n V_hig
+ 672.800001n V_hig
+ 672.900000n V_hig
+ 672.900001n V_hig
+ 673.000000n V_hig
+ 673.000001n V_hig
+ 673.100000n V_hig
+ 673.100001n V_hig
+ 673.200000n V_hig
+ 673.200001n V_hig
+ 673.300000n V_hig
+ 673.300001n V_hig
+ 673.400000n V_hig
+ 673.400001n V_hig
+ 673.500000n V_hig
+ 673.500001n V_hig
+ 673.600000n V_hig
+ 673.600001n V_hig
+ 673.700000n V_hig
+ 673.700001n V_hig
+ 673.800000n V_hig
+ 673.800001n V_hig
+ 673.900000n V_hig
+ 673.900001n V_hig
+ 674.000000n V_hig
+ 674.000001n V_hig
+ 674.100000n V_hig
+ 674.100001n V_hig
+ 674.200000n V_hig
+ 674.200001n V_hig
+ 674.300000n V_hig
+ 674.300001n V_hig
+ 674.400000n V_hig
+ 674.400001n V_hig
+ 674.500000n V_hig
+ 674.500001n V_hig
+ 674.600000n V_hig
+ 674.600001n V_hig
+ 674.700000n V_hig
+ 674.700001n V_hig
+ 674.800000n V_hig
+ 674.800001n V_hig
+ 674.900000n V_hig
+ 674.900001n V_hig
+ 675.000000n V_hig
+ 675.000001n V_low
+ 675.100000n V_low
+ 675.100001n V_low
+ 675.200000n V_low
+ 675.200001n V_low
+ 675.300000n V_low
+ 675.300001n V_low
+ 675.400000n V_low
+ 675.400001n V_low
+ 675.500000n V_low
+ 675.500001n V_low
+ 675.600000n V_low
+ 675.600001n V_low
+ 675.700000n V_low
+ 675.700001n V_low
+ 675.800000n V_low
+ 675.800001n V_low
+ 675.900000n V_low
+ 675.900001n V_low
+ 676.000000n V_low
+ 676.000001n V_low
+ 676.100000n V_low
+ 676.100001n V_low
+ 676.200000n V_low
+ 676.200001n V_low
+ 676.300000n V_low
+ 676.300001n V_low
+ 676.400000n V_low
+ 676.400001n V_low
+ 676.500000n V_low
+ 676.500001n V_low
+ 676.600000n V_low
+ 676.600001n V_low
+ 676.700000n V_low
+ 676.700001n V_low
+ 676.800000n V_low
+ 676.800001n V_low
+ 676.900000n V_low
+ 676.900001n V_low
+ 677.000000n V_low
+ 677.000001n V_hig
+ 677.100000n V_hig
+ 677.100001n V_hig
+ 677.200000n V_hig
+ 677.200001n V_hig
+ 677.300000n V_hig
+ 677.300001n V_hig
+ 677.400000n V_hig
+ 677.400001n V_hig
+ 677.500000n V_hig
+ 677.500001n V_hig
+ 677.600000n V_hig
+ 677.600001n V_hig
+ 677.700000n V_hig
+ 677.700001n V_hig
+ 677.800000n V_hig
+ 677.800001n V_hig
+ 677.900000n V_hig
+ 677.900001n V_hig
+ 678.000000n V_hig
+ 678.000001n V_low
+ 678.100000n V_low
+ 678.100001n V_low
+ 678.200000n V_low
+ 678.200001n V_low
+ 678.300000n V_low
+ 678.300001n V_low
+ 678.400000n V_low
+ 678.400001n V_low
+ 678.500000n V_low
+ 678.500001n V_low
+ 678.600000n V_low
+ 678.600001n V_low
+ 678.700000n V_low
+ 678.700001n V_low
+ 678.800000n V_low
+ 678.800001n V_low
+ 678.900000n V_low
+ 678.900001n V_low
+ 679.000000n V_low
+ 679.000001n V_hig
+ 679.100000n V_hig
+ 679.100001n V_hig
+ 679.200000n V_hig
+ 679.200001n V_hig
+ 679.300000n V_hig
+ 679.300001n V_hig
+ 679.400000n V_hig
+ 679.400001n V_hig
+ 679.500000n V_hig
+ 679.500001n V_hig
+ 679.600000n V_hig
+ 679.600001n V_hig
+ 679.700000n V_hig
+ 679.700001n V_hig
+ 679.800000n V_hig
+ 679.800001n V_hig
+ 679.900000n V_hig
+ 679.900001n V_hig
+ 680.000000n V_hig
+ 680.000001n V_low
+ 680.100000n V_low
+ 680.100001n V_low
+ 680.200000n V_low
+ 680.200001n V_low
+ 680.300000n V_low
+ 680.300001n V_low
+ 680.400000n V_low
+ 680.400001n V_low
+ 680.500000n V_low
+ 680.500001n V_low
+ 680.600000n V_low
+ 680.600001n V_low
+ 680.700000n V_low
+ 680.700001n V_low
+ 680.800000n V_low
+ 680.800001n V_low
+ 680.900000n V_low
+ 680.900001n V_low
+ 681.000000n V_low
+ 681.000001n V_hig
+ 681.100000n V_hig
+ 681.100001n V_hig
+ 681.200000n V_hig
+ 681.200001n V_hig
+ 681.300000n V_hig
+ 681.300001n V_hig
+ 681.400000n V_hig
+ 681.400001n V_hig
+ 681.500000n V_hig
+ 681.500001n V_hig
+ 681.600000n V_hig
+ 681.600001n V_hig
+ 681.700000n V_hig
+ 681.700001n V_hig
+ 681.800000n V_hig
+ 681.800001n V_hig
+ 681.900000n V_hig
+ 681.900001n V_hig
+ 682.000000n V_hig
+ 682.000001n V_hig
+ 682.100000n V_hig
+ 682.100001n V_hig
+ 682.200000n V_hig
+ 682.200001n V_hig
+ 682.300000n V_hig
+ 682.300001n V_hig
+ 682.400000n V_hig
+ 682.400001n V_hig
+ 682.500000n V_hig
+ 682.500001n V_hig
+ 682.600000n V_hig
+ 682.600001n V_hig
+ 682.700000n V_hig
+ 682.700001n V_hig
+ 682.800000n V_hig
+ 682.800001n V_hig
+ 682.900000n V_hig
+ 682.900001n V_hig
+ 683.000000n V_hig
+ 683.000001n V_low
+ 683.100000n V_low
+ 683.100001n V_low
+ 683.200000n V_low
+ 683.200001n V_low
+ 683.300000n V_low
+ 683.300001n V_low
+ 683.400000n V_low
+ 683.400001n V_low
+ 683.500000n V_low
+ 683.500001n V_low
+ 683.600000n V_low
+ 683.600001n V_low
+ 683.700000n V_low
+ 683.700001n V_low
+ 683.800000n V_low
+ 683.800001n V_low
+ 683.900000n V_low
+ 683.900001n V_low
+ 684.000000n V_low
+ 684.000001n V_hig
+ 684.100000n V_hig
+ 684.100001n V_hig
+ 684.200000n V_hig
+ 684.200001n V_hig
+ 684.300000n V_hig
+ 684.300001n V_hig
+ 684.400000n V_hig
+ 684.400001n V_hig
+ 684.500000n V_hig
+ 684.500001n V_hig
+ 684.600000n V_hig
+ 684.600001n V_hig
+ 684.700000n V_hig
+ 684.700001n V_hig
+ 684.800000n V_hig
+ 684.800001n V_hig
+ 684.900000n V_hig
+ 684.900001n V_hig
+ 685.000000n V_hig
+ 685.000001n V_hig
+ 685.100000n V_hig
+ 685.100001n V_hig
+ 685.200000n V_hig
+ 685.200001n V_hig
+ 685.300000n V_hig
+ 685.300001n V_hig
+ 685.400000n V_hig
+ 685.400001n V_hig
+ 685.500000n V_hig
+ 685.500001n V_hig
+ 685.600000n V_hig
+ 685.600001n V_hig
+ 685.700000n V_hig
+ 685.700001n V_hig
+ 685.800000n V_hig
+ 685.800001n V_hig
+ 685.900000n V_hig
+ 685.900001n V_hig
+ 686.000000n V_hig
+ 686.000001n V_hig
+ 686.100000n V_hig
+ 686.100001n V_hig
+ 686.200000n V_hig
+ 686.200001n V_hig
+ 686.300000n V_hig
+ 686.300001n V_hig
+ 686.400000n V_hig
+ 686.400001n V_hig
+ 686.500000n V_hig
+ 686.500001n V_hig
+ 686.600000n V_hig
+ 686.600001n V_hig
+ 686.700000n V_hig
+ 686.700001n V_hig
+ 686.800000n V_hig
+ 686.800001n V_hig
+ 686.900000n V_hig
+ 686.900001n V_hig
+ 687.000000n V_hig
+ 687.000001n V_hig
+ 687.100000n V_hig
+ 687.100001n V_hig
+ 687.200000n V_hig
+ 687.200001n V_hig
+ 687.300000n V_hig
+ 687.300001n V_hig
+ 687.400000n V_hig
+ 687.400001n V_hig
+ 687.500000n V_hig
+ 687.500001n V_hig
+ 687.600000n V_hig
+ 687.600001n V_hig
+ 687.700000n V_hig
+ 687.700001n V_hig
+ 687.800000n V_hig
+ 687.800001n V_hig
+ 687.900000n V_hig
+ 687.900001n V_hig
+ 688.000000n V_hig
+ 688.000001n V_hig
+ 688.100000n V_hig
+ 688.100001n V_hig
+ 688.200000n V_hig
+ 688.200001n V_hig
+ 688.300000n V_hig
+ 688.300001n V_hig
+ 688.400000n V_hig
+ 688.400001n V_hig
+ 688.500000n V_hig
+ 688.500001n V_hig
+ 688.600000n V_hig
+ 688.600001n V_hig
+ 688.700000n V_hig
+ 688.700001n V_hig
+ 688.800000n V_hig
+ 688.800001n V_hig
+ 688.900000n V_hig
+ 688.900001n V_hig
+ 689.000000n V_hig
+ 689.000001n V_hig
+ 689.100000n V_hig
+ 689.100001n V_hig
+ 689.200000n V_hig
+ 689.200001n V_hig
+ 689.300000n V_hig
+ 689.300001n V_hig
+ 689.400000n V_hig
+ 689.400001n V_hig
+ 689.500000n V_hig
+ 689.500001n V_hig
+ 689.600000n V_hig
+ 689.600001n V_hig
+ 689.700000n V_hig
+ 689.700001n V_hig
+ 689.800000n V_hig
+ 689.800001n V_hig
+ 689.900000n V_hig
+ 689.900001n V_hig
+ 690.000000n V_hig
+ 690.000001n V_low
+ 690.100000n V_low
+ 690.100001n V_low
+ 690.200000n V_low
+ 690.200001n V_low
+ 690.300000n V_low
+ 690.300001n V_low
+ 690.400000n V_low
+ 690.400001n V_low
+ 690.500000n V_low
+ 690.500001n V_low
+ 690.600000n V_low
+ 690.600001n V_low
+ 690.700000n V_low
+ 690.700001n V_low
+ 690.800000n V_low
+ 690.800001n V_low
+ 690.900000n V_low
+ 690.900001n V_low
+ 691.000000n V_low
+ 691.000001n V_low
+ 691.100000n V_low
+ 691.100001n V_low
+ 691.200000n V_low
+ 691.200001n V_low
+ 691.300000n V_low
+ 691.300001n V_low
+ 691.400000n V_low
+ 691.400001n V_low
+ 691.500000n V_low
+ 691.500001n V_low
+ 691.600000n V_low
+ 691.600001n V_low
+ 691.700000n V_low
+ 691.700001n V_low
+ 691.800000n V_low
+ 691.800001n V_low
+ 691.900000n V_low
+ 691.900001n V_low
+ 692.000000n V_low
+ 692.000001n V_hig
+ 692.100000n V_hig
+ 692.100001n V_hig
+ 692.200000n V_hig
+ 692.200001n V_hig
+ 692.300000n V_hig
+ 692.300001n V_hig
+ 692.400000n V_hig
+ 692.400001n V_hig
+ 692.500000n V_hig
+ 692.500001n V_hig
+ 692.600000n V_hig
+ 692.600001n V_hig
+ 692.700000n V_hig
+ 692.700001n V_hig
+ 692.800000n V_hig
+ 692.800001n V_hig
+ 692.900000n V_hig
+ 692.900001n V_hig
+ 693.000000n V_hig
+ 693.000001n V_low
+ 693.100000n V_low
+ 693.100001n V_low
+ 693.200000n V_low
+ 693.200001n V_low
+ 693.300000n V_low
+ 693.300001n V_low
+ 693.400000n V_low
+ 693.400001n V_low
+ 693.500000n V_low
+ 693.500001n V_low
+ 693.600000n V_low
+ 693.600001n V_low
+ 693.700000n V_low
+ 693.700001n V_low
+ 693.800000n V_low
+ 693.800001n V_low
+ 693.900000n V_low
+ 693.900001n V_low
+ 694.000000n V_low
+ 694.000001n V_low
+ 694.100000n V_low
+ 694.100001n V_low
+ 694.200000n V_low
+ 694.200001n V_low
+ 694.300000n V_low
+ 694.300001n V_low
+ 694.400000n V_low
+ 694.400001n V_low
+ 694.500000n V_low
+ 694.500001n V_low
+ 694.600000n V_low
+ 694.600001n V_low
+ 694.700000n V_low
+ 694.700001n V_low
+ 694.800000n V_low
+ 694.800001n V_low
+ 694.900000n V_low
+ 694.900001n V_low
+ 695.000000n V_low
+ 695.000001n V_low
+ 695.100000n V_low
+ 695.100001n V_low
+ 695.200000n V_low
+ 695.200001n V_low
+ 695.300000n V_low
+ 695.300001n V_low
+ 695.400000n V_low
+ 695.400001n V_low
+ 695.500000n V_low
+ 695.500001n V_low
+ 695.600000n V_low
+ 695.600001n V_low
+ 695.700000n V_low
+ 695.700001n V_low
+ 695.800000n V_low
+ 695.800001n V_low
+ 695.900000n V_low
+ 695.900001n V_low
+ 696.000000n V_low
+ 696.000001n V_low
+ 696.100000n V_low
+ 696.100001n V_low
+ 696.200000n V_low
+ 696.200001n V_low
+ 696.300000n V_low
+ 696.300001n V_low
+ 696.400000n V_low
+ 696.400001n V_low
+ 696.500000n V_low
+ 696.500001n V_low
+ 696.600000n V_low
+ 696.600001n V_low
+ 696.700000n V_low
+ 696.700001n V_low
+ 696.800000n V_low
+ 696.800001n V_low
+ 696.900000n V_low
+ 696.900001n V_low
+ 697.000000n V_low
+ 697.000001n V_low
+ 697.100000n V_low
+ 697.100001n V_low
+ 697.200000n V_low
+ 697.200001n V_low
+ 697.300000n V_low
+ 697.300001n V_low
+ 697.400000n V_low
+ 697.400001n V_low
+ 697.500000n V_low
+ 697.500001n V_low
+ 697.600000n V_low
+ 697.600001n V_low
+ 697.700000n V_low
+ 697.700001n V_low
+ 697.800000n V_low
+ 697.800001n V_low
+ 697.900000n V_low
+ 697.900001n V_low
+ 698.000000n V_low
+ 698.000001n V_low
+ 698.100000n V_low
+ 698.100001n V_low
+ 698.200000n V_low
+ 698.200001n V_low
+ 698.300000n V_low
+ 698.300001n V_low
+ 698.400000n V_low
+ 698.400001n V_low
+ 698.500000n V_low
+ 698.500001n V_low
+ 698.600000n V_low
+ 698.600001n V_low
+ 698.700000n V_low
+ 698.700001n V_low
+ 698.800000n V_low
+ 698.800001n V_low
+ 698.900000n V_low
+ 698.900001n V_low
+ 699.000000n V_low
+ 699.000001n V_hig
+ 699.100000n V_hig
+ 699.100001n V_hig
+ 699.200000n V_hig
+ 699.200001n V_hig
+ 699.300000n V_hig
+ 699.300001n V_hig
+ 699.400000n V_hig
+ 699.400001n V_hig
+ 699.500000n V_hig
+ 699.500001n V_hig
+ 699.600000n V_hig
+ 699.600001n V_hig
+ 699.700000n V_hig
+ 699.700001n V_hig
+ 699.800000n V_hig
+ 699.800001n V_hig
+ 699.900000n V_hig
+ 699.900001n V_hig
+ 700.000000n V_hig
+ 700.000001n V_low
+ 700.100000n V_low
+ 700.100001n V_low
+ 700.200000n V_low
+ 700.200001n V_low
+ 700.300000n V_low
+ 700.300001n V_low
+ 700.400000n V_low
+ 700.400001n V_low
+ 700.500000n V_low
+ 700.500001n V_low
+ 700.600000n V_low
+ 700.600001n V_low
+ 700.700000n V_low
+ 700.700001n V_low
+ 700.800000n V_low
+ 700.800001n V_low
+ 700.900000n V_low
+ 700.900001n V_low
+ 701.000000n V_low
+ 701.000001n V_low
+ 701.100000n V_low
+ 701.100001n V_low
+ 701.200000n V_low
+ 701.200001n V_low
+ 701.300000n V_low
+ 701.300001n V_low
+ 701.400000n V_low
+ 701.400001n V_low
+ 701.500000n V_low
+ 701.500001n V_low
+ 701.600000n V_low
+ 701.600001n V_low
+ 701.700000n V_low
+ 701.700001n V_low
+ 701.800000n V_low
+ 701.800001n V_low
+ 701.900000n V_low
+ 701.900001n V_low
+ 702.000000n V_low
+ 702.000001n V_low
+ 702.100000n V_low
+ 702.100001n V_low
+ 702.200000n V_low
+ 702.200001n V_low
+ 702.300000n V_low
+ 702.300001n V_low
+ 702.400000n V_low
+ 702.400001n V_low
+ 702.500000n V_low
+ 702.500001n V_low
+ 702.600000n V_low
+ 702.600001n V_low
+ 702.700000n V_low
+ 702.700001n V_low
+ 702.800000n V_low
+ 702.800001n V_low
+ 702.900000n V_low
+ 702.900001n V_low
+ 703.000000n V_low
+ 703.000001n V_hig
+ 703.100000n V_hig
+ 703.100001n V_hig
+ 703.200000n V_hig
+ 703.200001n V_hig
+ 703.300000n V_hig
+ 703.300001n V_hig
+ 703.400000n V_hig
+ 703.400001n V_hig
+ 703.500000n V_hig
+ 703.500001n V_hig
+ 703.600000n V_hig
+ 703.600001n V_hig
+ 703.700000n V_hig
+ 703.700001n V_hig
+ 703.800000n V_hig
+ 703.800001n V_hig
+ 703.900000n V_hig
+ 703.900001n V_hig
+ 704.000000n V_hig
+ 704.000001n V_low
+ 704.100000n V_low
+ 704.100001n V_low
+ 704.200000n V_low
+ 704.200001n V_low
+ 704.300000n V_low
+ 704.300001n V_low
+ 704.400000n V_low
+ 704.400001n V_low
+ 704.500000n V_low
+ 704.500001n V_low
+ 704.600000n V_low
+ 704.600001n V_low
+ 704.700000n V_low
+ 704.700001n V_low
+ 704.800000n V_low
+ 704.800001n V_low
+ 704.900000n V_low
+ 704.900001n V_low
+ 705.000000n V_low
+ 705.000001n V_low
+ 705.100000n V_low
+ 705.100001n V_low
+ 705.200000n V_low
+ 705.200001n V_low
+ 705.300000n V_low
+ 705.300001n V_low
+ 705.400000n V_low
+ 705.400001n V_low
+ 705.500000n V_low
+ 705.500001n V_low
+ 705.600000n V_low
+ 705.600001n V_low
+ 705.700000n V_low
+ 705.700001n V_low
+ 705.800000n V_low
+ 705.800001n V_low
+ 705.900000n V_low
+ 705.900001n V_low
+ 706.000000n V_low
+ 706.000001n V_low
+ 706.100000n V_low
+ 706.100001n V_low
+ 706.200000n V_low
+ 706.200001n V_low
+ 706.300000n V_low
+ 706.300001n V_low
+ 706.400000n V_low
+ 706.400001n V_low
+ 706.500000n V_low
+ 706.500001n V_low
+ 706.600000n V_low
+ 706.600001n V_low
+ 706.700000n V_low
+ 706.700001n V_low
+ 706.800000n V_low
+ 706.800001n V_low
+ 706.900000n V_low
+ 706.900001n V_low
+ 707.000000n V_low
+ 707.000001n V_low
+ 707.100000n V_low
+ 707.100001n V_low
+ 707.200000n V_low
+ 707.200001n V_low
+ 707.300000n V_low
+ 707.300001n V_low
+ 707.400000n V_low
+ 707.400001n V_low
+ 707.500000n V_low
+ 707.500001n V_low
+ 707.600000n V_low
+ 707.600001n V_low
+ 707.700000n V_low
+ 707.700001n V_low
+ 707.800000n V_low
+ 707.800001n V_low
+ 707.900000n V_low
+ 707.900001n V_low
+ 708.000000n V_low
+ 708.000001n V_hig
+ 708.100000n V_hig
+ 708.100001n V_hig
+ 708.200000n V_hig
+ 708.200001n V_hig
+ 708.300000n V_hig
+ 708.300001n V_hig
+ 708.400000n V_hig
+ 708.400001n V_hig
+ 708.500000n V_hig
+ 708.500001n V_hig
+ 708.600000n V_hig
+ 708.600001n V_hig
+ 708.700000n V_hig
+ 708.700001n V_hig
+ 708.800000n V_hig
+ 708.800001n V_hig
+ 708.900000n V_hig
+ 708.900001n V_hig
+ 709.000000n V_hig
+ 709.000001n V_hig
+ 709.100000n V_hig
+ 709.100001n V_hig
+ 709.200000n V_hig
+ 709.200001n V_hig
+ 709.300000n V_hig
+ 709.300001n V_hig
+ 709.400000n V_hig
+ 709.400001n V_hig
+ 709.500000n V_hig
+ 709.500001n V_hig
+ 709.600000n V_hig
+ 709.600001n V_hig
+ 709.700000n V_hig
+ 709.700001n V_hig
+ 709.800000n V_hig
+ 709.800001n V_hig
+ 709.900000n V_hig
+ 709.900001n V_hig
+ 710.000000n V_hig
+ 710.000001n V_low
+ 710.100000n V_low
+ 710.100001n V_low
+ 710.200000n V_low
+ 710.200001n V_low
+ 710.300000n V_low
+ 710.300001n V_low
+ 710.400000n V_low
+ 710.400001n V_low
+ 710.500000n V_low
+ 710.500001n V_low
+ 710.600000n V_low
+ 710.600001n V_low
+ 710.700000n V_low
+ 710.700001n V_low
+ 710.800000n V_low
+ 710.800001n V_low
+ 710.900000n V_low
+ 710.900001n V_low
+ 711.000000n V_low
+ 711.000001n V_low
+ 711.100000n V_low
+ 711.100001n V_low
+ 711.200000n V_low
+ 711.200001n V_low
+ 711.300000n V_low
+ 711.300001n V_low
+ 711.400000n V_low
+ 711.400001n V_low
+ 711.500000n V_low
+ 711.500001n V_low
+ 711.600000n V_low
+ 711.600001n V_low
+ 711.700000n V_low
+ 711.700001n V_low
+ 711.800000n V_low
+ 711.800001n V_low
+ 711.900000n V_low
+ 711.900001n V_low
+ 712.000000n V_low
+ 712.000001n V_low
+ 712.100000n V_low
+ 712.100001n V_low
+ 712.200000n V_low
+ 712.200001n V_low
+ 712.300000n V_low
+ 712.300001n V_low
+ 712.400000n V_low
+ 712.400001n V_low
+ 712.500000n V_low
+ 712.500001n V_low
+ 712.600000n V_low
+ 712.600001n V_low
+ 712.700000n V_low
+ 712.700001n V_low
+ 712.800000n V_low
+ 712.800001n V_low
+ 712.900000n V_low
+ 712.900001n V_low
+ 713.000000n V_low
+ 713.000001n V_low
+ 713.100000n V_low
+ 713.100001n V_low
+ 713.200000n V_low
+ 713.200001n V_low
+ 713.300000n V_low
+ 713.300001n V_low
+ 713.400000n V_low
+ 713.400001n V_low
+ 713.500000n V_low
+ 713.500001n V_low
+ 713.600000n V_low
+ 713.600001n V_low
+ 713.700000n V_low
+ 713.700001n V_low
+ 713.800000n V_low
+ 713.800001n V_low
+ 713.900000n V_low
+ 713.900001n V_low
+ 714.000000n V_low
+ 714.000001n V_hig
+ 714.100000n V_hig
+ 714.100001n V_hig
+ 714.200000n V_hig
+ 714.200001n V_hig
+ 714.300000n V_hig
+ 714.300001n V_hig
+ 714.400000n V_hig
+ 714.400001n V_hig
+ 714.500000n V_hig
+ 714.500001n V_hig
+ 714.600000n V_hig
+ 714.600001n V_hig
+ 714.700000n V_hig
+ 714.700001n V_hig
+ 714.800000n V_hig
+ 714.800001n V_hig
+ 714.900000n V_hig
+ 714.900001n V_hig
+ 715.000000n V_hig
+ 715.000001n V_hig
+ 715.100000n V_hig
+ 715.100001n V_hig
+ 715.200000n V_hig
+ 715.200001n V_hig
+ 715.300000n V_hig
+ 715.300001n V_hig
+ 715.400000n V_hig
+ 715.400001n V_hig
+ 715.500000n V_hig
+ 715.500001n V_hig
+ 715.600000n V_hig
+ 715.600001n V_hig
+ 715.700000n V_hig
+ 715.700001n V_hig
+ 715.800000n V_hig
+ 715.800001n V_hig
+ 715.900000n V_hig
+ 715.900001n V_hig
+ 716.000000n V_hig
+ 716.000001n V_hig
+ 716.100000n V_hig
+ 716.100001n V_hig
+ 716.200000n V_hig
+ 716.200001n V_hig
+ 716.300000n V_hig
+ 716.300001n V_hig
+ 716.400000n V_hig
+ 716.400001n V_hig
+ 716.500000n V_hig
+ 716.500001n V_hig
+ 716.600000n V_hig
+ 716.600001n V_hig
+ 716.700000n V_hig
+ 716.700001n V_hig
+ 716.800000n V_hig
+ 716.800001n V_hig
+ 716.900000n V_hig
+ 716.900001n V_hig
+ 717.000000n V_hig
+ 717.000001n V_hig
+ 717.100000n V_hig
+ 717.100001n V_hig
+ 717.200000n V_hig
+ 717.200001n V_hig
+ 717.300000n V_hig
+ 717.300001n V_hig
+ 717.400000n V_hig
+ 717.400001n V_hig
+ 717.500000n V_hig
+ 717.500001n V_hig
+ 717.600000n V_hig
+ 717.600001n V_hig
+ 717.700000n V_hig
+ 717.700001n V_hig
+ 717.800000n V_hig
+ 717.800001n V_hig
+ 717.900000n V_hig
+ 717.900001n V_hig
+ 718.000000n V_hig
+ 718.000001n V_low
+ 718.100000n V_low
+ 718.100001n V_low
+ 718.200000n V_low
+ 718.200001n V_low
+ 718.300000n V_low
+ 718.300001n V_low
+ 718.400000n V_low
+ 718.400001n V_low
+ 718.500000n V_low
+ 718.500001n V_low
+ 718.600000n V_low
+ 718.600001n V_low
+ 718.700000n V_low
+ 718.700001n V_low
+ 718.800000n V_low
+ 718.800001n V_low
+ 718.900000n V_low
+ 718.900001n V_low
+ 719.000000n V_low
+ 719.000001n V_low
+ 719.100000n V_low
+ 719.100001n V_low
+ 719.200000n V_low
+ 719.200001n V_low
+ 719.300000n V_low
+ 719.300001n V_low
+ 719.400000n V_low
+ 719.400001n V_low
+ 719.500000n V_low
+ 719.500001n V_low
+ 719.600000n V_low
+ 719.600001n V_low
+ 719.700000n V_low
+ 719.700001n V_low
+ 719.800000n V_low
+ 719.800001n V_low
+ 719.900000n V_low
+ 719.900001n V_low
+ 720.000000n V_low
+ 720.000001n V_low
+ 720.100000n V_low
+ 720.100001n V_low
+ 720.200000n V_low
+ 720.200001n V_low
+ 720.300000n V_low
+ 720.300001n V_low
+ 720.400000n V_low
+ 720.400001n V_low
+ 720.500000n V_low
+ 720.500001n V_low
+ 720.600000n V_low
+ 720.600001n V_low
+ 720.700000n V_low
+ 720.700001n V_low
+ 720.800000n V_low
+ 720.800001n V_low
+ 720.900000n V_low
+ 720.900001n V_low
+ 721.000000n V_low
+ 721.000001n V_hig
+ 721.100000n V_hig
+ 721.100001n V_hig
+ 721.200000n V_hig
+ 721.200001n V_hig
+ 721.300000n V_hig
+ 721.300001n V_hig
+ 721.400000n V_hig
+ 721.400001n V_hig
+ 721.500000n V_hig
+ 721.500001n V_hig
+ 721.600000n V_hig
+ 721.600001n V_hig
+ 721.700000n V_hig
+ 721.700001n V_hig
+ 721.800000n V_hig
+ 721.800001n V_hig
+ 721.900000n V_hig
+ 721.900001n V_hig
+ 722.000000n V_hig
+ 722.000001n V_low
+ 722.100000n V_low
+ 722.100001n V_low
+ 722.200000n V_low
+ 722.200001n V_low
+ 722.300000n V_low
+ 722.300001n V_low
+ 722.400000n V_low
+ 722.400001n V_low
+ 722.500000n V_low
+ 722.500001n V_low
+ 722.600000n V_low
+ 722.600001n V_low
+ 722.700000n V_low
+ 722.700001n V_low
+ 722.800000n V_low
+ 722.800001n V_low
+ 722.900000n V_low
+ 722.900001n V_low
+ 723.000000n V_low
+ 723.000001n V_low
+ 723.100000n V_low
+ 723.100001n V_low
+ 723.200000n V_low
+ 723.200001n V_low
+ 723.300000n V_low
+ 723.300001n V_low
+ 723.400000n V_low
+ 723.400001n V_low
+ 723.500000n V_low
+ 723.500001n V_low
+ 723.600000n V_low
+ 723.600001n V_low
+ 723.700000n V_low
+ 723.700001n V_low
+ 723.800000n V_low
+ 723.800001n V_low
+ 723.900000n V_low
+ 723.900001n V_low
+ 724.000000n V_low
+ 724.000001n V_hig
+ 724.100000n V_hig
+ 724.100001n V_hig
+ 724.200000n V_hig
+ 724.200001n V_hig
+ 724.300000n V_hig
+ 724.300001n V_hig
+ 724.400000n V_hig
+ 724.400001n V_hig
+ 724.500000n V_hig
+ 724.500001n V_hig
+ 724.600000n V_hig
+ 724.600001n V_hig
+ 724.700000n V_hig
+ 724.700001n V_hig
+ 724.800000n V_hig
+ 724.800001n V_hig
+ 724.900000n V_hig
+ 724.900001n V_hig
+ 725.000000n V_hig
+ 725.000001n V_hig
+ 725.100000n V_hig
+ 725.100001n V_hig
+ 725.200000n V_hig
+ 725.200001n V_hig
+ 725.300000n V_hig
+ 725.300001n V_hig
+ 725.400000n V_hig
+ 725.400001n V_hig
+ 725.500000n V_hig
+ 725.500001n V_hig
+ 725.600000n V_hig
+ 725.600001n V_hig
+ 725.700000n V_hig
+ 725.700001n V_hig
+ 725.800000n V_hig
+ 725.800001n V_hig
+ 725.900000n V_hig
+ 725.900001n V_hig
+ 726.000000n V_hig
+ 726.000001n V_hig
+ 726.100000n V_hig
+ 726.100001n V_hig
+ 726.200000n V_hig
+ 726.200001n V_hig
+ 726.300000n V_hig
+ 726.300001n V_hig
+ 726.400000n V_hig
+ 726.400001n V_hig
+ 726.500000n V_hig
+ 726.500001n V_hig
+ 726.600000n V_hig
+ 726.600001n V_hig
+ 726.700000n V_hig
+ 726.700001n V_hig
+ 726.800000n V_hig
+ 726.800001n V_hig
+ 726.900000n V_hig
+ 726.900001n V_hig
+ 727.000000n V_hig
+ 727.000001n V_hig
+ 727.100000n V_hig
+ 727.100001n V_hig
+ 727.200000n V_hig
+ 727.200001n V_hig
+ 727.300000n V_hig
+ 727.300001n V_hig
+ 727.400000n V_hig
+ 727.400001n V_hig
+ 727.500000n V_hig
+ 727.500001n V_hig
+ 727.600000n V_hig
+ 727.600001n V_hig
+ 727.700000n V_hig
+ 727.700001n V_hig
+ 727.800000n V_hig
+ 727.800001n V_hig
+ 727.900000n V_hig
+ 727.900001n V_hig
+ 728.000000n V_hig
+ 728.000001n V_low
+ 728.100000n V_low
+ 728.100001n V_low
+ 728.200000n V_low
+ 728.200001n V_low
+ 728.300000n V_low
+ 728.300001n V_low
+ 728.400000n V_low
+ 728.400001n V_low
+ 728.500000n V_low
+ 728.500001n V_low
+ 728.600000n V_low
+ 728.600001n V_low
+ 728.700000n V_low
+ 728.700001n V_low
+ 728.800000n V_low
+ 728.800001n V_low
+ 728.900000n V_low
+ 728.900001n V_low
+ 729.000000n V_low
+ 729.000001n V_hig
+ 729.100000n V_hig
+ 729.100001n V_hig
+ 729.200000n V_hig
+ 729.200001n V_hig
+ 729.300000n V_hig
+ 729.300001n V_hig
+ 729.400000n V_hig
+ 729.400001n V_hig
+ 729.500000n V_hig
+ 729.500001n V_hig
+ 729.600000n V_hig
+ 729.600001n V_hig
+ 729.700000n V_hig
+ 729.700001n V_hig
+ 729.800000n V_hig
+ 729.800001n V_hig
+ 729.900000n V_hig
+ 729.900001n V_hig
+ 730.000000n V_hig
+ 730.000001n V_hig
+ 730.100000n V_hig
+ 730.100001n V_hig
+ 730.200000n V_hig
+ 730.200001n V_hig
+ 730.300000n V_hig
+ 730.300001n V_hig
+ 730.400000n V_hig
+ 730.400001n V_hig
+ 730.500000n V_hig
+ 730.500001n V_hig
+ 730.600000n V_hig
+ 730.600001n V_hig
+ 730.700000n V_hig
+ 730.700001n V_hig
+ 730.800000n V_hig
+ 730.800001n V_hig
+ 730.900000n V_hig
+ 730.900001n V_hig
+ 731.000000n V_hig
+ 731.000001n V_low
+ 731.100000n V_low
+ 731.100001n V_low
+ 731.200000n V_low
+ 731.200001n V_low
+ 731.300000n V_low
+ 731.300001n V_low
+ 731.400000n V_low
+ 731.400001n V_low
+ 731.500000n V_low
+ 731.500001n V_low
+ 731.600000n V_low
+ 731.600001n V_low
+ 731.700000n V_low
+ 731.700001n V_low
+ 731.800000n V_low
+ 731.800001n V_low
+ 731.900000n V_low
+ 731.900001n V_low
+ 732.000000n V_low
+ 732.000001n V_low
+ 732.100000n V_low
+ 732.100001n V_low
+ 732.200000n V_low
+ 732.200001n V_low
+ 732.300000n V_low
+ 732.300001n V_low
+ 732.400000n V_low
+ 732.400001n V_low
+ 732.500000n V_low
+ 732.500001n V_low
+ 732.600000n V_low
+ 732.600001n V_low
+ 732.700000n V_low
+ 732.700001n V_low
+ 732.800000n V_low
+ 732.800001n V_low
+ 732.900000n V_low
+ 732.900001n V_low
+ 733.000000n V_low
+ 733.000001n V_hig
+ 733.100000n V_hig
+ 733.100001n V_hig
+ 733.200000n V_hig
+ 733.200001n V_hig
+ 733.300000n V_hig
+ 733.300001n V_hig
+ 733.400000n V_hig
+ 733.400001n V_hig
+ 733.500000n V_hig
+ 733.500001n V_hig
+ 733.600000n V_hig
+ 733.600001n V_hig
+ 733.700000n V_hig
+ 733.700001n V_hig
+ 733.800000n V_hig
+ 733.800001n V_hig
+ 733.900000n V_hig
+ 733.900001n V_hig
+ 734.000000n V_hig
+ 734.000001n V_hig
+ 734.100000n V_hig
+ 734.100001n V_hig
+ 734.200000n V_hig
+ 734.200001n V_hig
+ 734.300000n V_hig
+ 734.300001n V_hig
+ 734.400000n V_hig
+ 734.400001n V_hig
+ 734.500000n V_hig
+ 734.500001n V_hig
+ 734.600000n V_hig
+ 734.600001n V_hig
+ 734.700000n V_hig
+ 734.700001n V_hig
+ 734.800000n V_hig
+ 734.800001n V_hig
+ 734.900000n V_hig
+ 734.900001n V_hig
+ 735.000000n V_hig
+ 735.000001n V_low
+ 735.100000n V_low
+ 735.100001n V_low
+ 735.200000n V_low
+ 735.200001n V_low
+ 735.300000n V_low
+ 735.300001n V_low
+ 735.400000n V_low
+ 735.400001n V_low
+ 735.500000n V_low
+ 735.500001n V_low
+ 735.600000n V_low
+ 735.600001n V_low
+ 735.700000n V_low
+ 735.700001n V_low
+ 735.800000n V_low
+ 735.800001n V_low
+ 735.900000n V_low
+ 735.900001n V_low
+ 736.000000n V_low
+ 736.000001n V_low
+ 736.100000n V_low
+ 736.100001n V_low
+ 736.200000n V_low
+ 736.200001n V_low
+ 736.300000n V_low
+ 736.300001n V_low
+ 736.400000n V_low
+ 736.400001n V_low
+ 736.500000n V_low
+ 736.500001n V_low
+ 736.600000n V_low
+ 736.600001n V_low
+ 736.700000n V_low
+ 736.700001n V_low
+ 736.800000n V_low
+ 736.800001n V_low
+ 736.900000n V_low
+ 736.900001n V_low
+ 737.000000n V_low
+ 737.000001n V_hig
+ 737.100000n V_hig
+ 737.100001n V_hig
+ 737.200000n V_hig
+ 737.200001n V_hig
+ 737.300000n V_hig
+ 737.300001n V_hig
+ 737.400000n V_hig
+ 737.400001n V_hig
+ 737.500000n V_hig
+ 737.500001n V_hig
+ 737.600000n V_hig
+ 737.600001n V_hig
+ 737.700000n V_hig
+ 737.700001n V_hig
+ 737.800000n V_hig
+ 737.800001n V_hig
+ 737.900000n V_hig
+ 737.900001n V_hig
+ 738.000000n V_hig
+ 738.000001n V_hig
+ 738.100000n V_hig
+ 738.100001n V_hig
+ 738.200000n V_hig
+ 738.200001n V_hig
+ 738.300000n V_hig
+ 738.300001n V_hig
+ 738.400000n V_hig
+ 738.400001n V_hig
+ 738.500000n V_hig
+ 738.500001n V_hig
+ 738.600000n V_hig
+ 738.600001n V_hig
+ 738.700000n V_hig
+ 738.700001n V_hig
+ 738.800000n V_hig
+ 738.800001n V_hig
+ 738.900000n V_hig
+ 738.900001n V_hig
+ 739.000000n V_hig
+ 739.000001n V_hig
+ 739.100000n V_hig
+ 739.100001n V_hig
+ 739.200000n V_hig
+ 739.200001n V_hig
+ 739.300000n V_hig
+ 739.300001n V_hig
+ 739.400000n V_hig
+ 739.400001n V_hig
+ 739.500000n V_hig
+ 739.500001n V_hig
+ 739.600000n V_hig
+ 739.600001n V_hig
+ 739.700000n V_hig
+ 739.700001n V_hig
+ 739.800000n V_hig
+ 739.800001n V_hig
+ 739.900000n V_hig
+ 739.900001n V_hig
+ 740.000000n V_hig
+ 740.000001n V_low
+ 740.100000n V_low
+ 740.100001n V_low
+ 740.200000n V_low
+ 740.200001n V_low
+ 740.300000n V_low
+ 740.300001n V_low
+ 740.400000n V_low
+ 740.400001n V_low
+ 740.500000n V_low
+ 740.500001n V_low
+ 740.600000n V_low
+ 740.600001n V_low
+ 740.700000n V_low
+ 740.700001n V_low
+ 740.800000n V_low
+ 740.800001n V_low
+ 740.900000n V_low
+ 740.900001n V_low
+ 741.000000n V_low
+ 741.000001n V_low
+ 741.100000n V_low
+ 741.100001n V_low
+ 741.200000n V_low
+ 741.200001n V_low
+ 741.300000n V_low
+ 741.300001n V_low
+ 741.400000n V_low
+ 741.400001n V_low
+ 741.500000n V_low
+ 741.500001n V_low
+ 741.600000n V_low
+ 741.600001n V_low
+ 741.700000n V_low
+ 741.700001n V_low
+ 741.800000n V_low
+ 741.800001n V_low
+ 741.900000n V_low
+ 741.900001n V_low
+ 742.000000n V_low
+ 742.000001n V_hig
+ 742.100000n V_hig
+ 742.100001n V_hig
+ 742.200000n V_hig
+ 742.200001n V_hig
+ 742.300000n V_hig
+ 742.300001n V_hig
+ 742.400000n V_hig
+ 742.400001n V_hig
+ 742.500000n V_hig
+ 742.500001n V_hig
+ 742.600000n V_hig
+ 742.600001n V_hig
+ 742.700000n V_hig
+ 742.700001n V_hig
+ 742.800000n V_hig
+ 742.800001n V_hig
+ 742.900000n V_hig
+ 742.900001n V_hig
+ 743.000000n V_hig
+ 743.000001n V_hig
+ 743.100000n V_hig
+ 743.100001n V_hig
+ 743.200000n V_hig
+ 743.200001n V_hig
+ 743.300000n V_hig
+ 743.300001n V_hig
+ 743.400000n V_hig
+ 743.400001n V_hig
+ 743.500000n V_hig
+ 743.500001n V_hig
+ 743.600000n V_hig
+ 743.600001n V_hig
+ 743.700000n V_hig
+ 743.700001n V_hig
+ 743.800000n V_hig
+ 743.800001n V_hig
+ 743.900000n V_hig
+ 743.900001n V_hig
+ 744.000000n V_hig
+ 744.000001n V_low
+ 744.100000n V_low
+ 744.100001n V_low
+ 744.200000n V_low
+ 744.200001n V_low
+ 744.300000n V_low
+ 744.300001n V_low
+ 744.400000n V_low
+ 744.400001n V_low
+ 744.500000n V_low
+ 744.500001n V_low
+ 744.600000n V_low
+ 744.600001n V_low
+ 744.700000n V_low
+ 744.700001n V_low
+ 744.800000n V_low
+ 744.800001n V_low
+ 744.900000n V_low
+ 744.900001n V_low
+ 745.000000n V_low
+ 745.000001n V_low
+ 745.100000n V_low
+ 745.100001n V_low
+ 745.200000n V_low
+ 745.200001n V_low
+ 745.300000n V_low
+ 745.300001n V_low
+ 745.400000n V_low
+ 745.400001n V_low
+ 745.500000n V_low
+ 745.500001n V_low
+ 745.600000n V_low
+ 745.600001n V_low
+ 745.700000n V_low
+ 745.700001n V_low
+ 745.800000n V_low
+ 745.800001n V_low
+ 745.900000n V_low
+ 745.900001n V_low
+ 746.000000n V_low
+ 746.000001n V_low
+ 746.100000n V_low
+ 746.100001n V_low
+ 746.200000n V_low
+ 746.200001n V_low
+ 746.300000n V_low
+ 746.300001n V_low
+ 746.400000n V_low
+ 746.400001n V_low
+ 746.500000n V_low
+ 746.500001n V_low
+ 746.600000n V_low
+ 746.600001n V_low
+ 746.700000n V_low
+ 746.700001n V_low
+ 746.800000n V_low
+ 746.800001n V_low
+ 746.900000n V_low
+ 746.900001n V_low
+ 747.000000n V_low
+ 747.000001n V_low
+ 747.100000n V_low
+ 747.100001n V_low
+ 747.200000n V_low
+ 747.200001n V_low
+ 747.300000n V_low
+ 747.300001n V_low
+ 747.400000n V_low
+ 747.400001n V_low
+ 747.500000n V_low
+ 747.500001n V_low
+ 747.600000n V_low
+ 747.600001n V_low
+ 747.700000n V_low
+ 747.700001n V_low
+ 747.800000n V_low
+ 747.800001n V_low
+ 747.900000n V_low
+ 747.900001n V_low
+ 748.000000n V_low
+ 748.000001n V_hig
+ 748.100000n V_hig
+ 748.100001n V_hig
+ 748.200000n V_hig
+ 748.200001n V_hig
+ 748.300000n V_hig
+ 748.300001n V_hig
+ 748.400000n V_hig
+ 748.400001n V_hig
+ 748.500000n V_hig
+ 748.500001n V_hig
+ 748.600000n V_hig
+ 748.600001n V_hig
+ 748.700000n V_hig
+ 748.700001n V_hig
+ 748.800000n V_hig
+ 748.800001n V_hig
+ 748.900000n V_hig
+ 748.900001n V_hig
+ 749.000000n V_hig
+ 749.000001n V_hig
+ 749.100000n V_hig
+ 749.100001n V_hig
+ 749.200000n V_hig
+ 749.200001n V_hig
+ 749.300000n V_hig
+ 749.300001n V_hig
+ 749.400000n V_hig
+ 749.400001n V_hig
+ 749.500000n V_hig
+ 749.500001n V_hig
+ 749.600000n V_hig
+ 749.600001n V_hig
+ 749.700000n V_hig
+ 749.700001n V_hig
+ 749.800000n V_hig
+ 749.800001n V_hig
+ 749.900000n V_hig
+ 749.900001n V_hig
+ 750.000000n V_hig
+ 750.000001n V_low
+ 750.100000n V_low
+ 750.100001n V_low
+ 750.200000n V_low
+ 750.200001n V_low
+ 750.300000n V_low
+ 750.300001n V_low
+ 750.400000n V_low
+ 750.400001n V_low
+ 750.500000n V_low
+ 750.500001n V_low
+ 750.600000n V_low
+ 750.600001n V_low
+ 750.700000n V_low
+ 750.700001n V_low
+ 750.800000n V_low
+ 750.800001n V_low
+ 750.900000n V_low
+ 750.900001n V_low
+ 751.000000n V_low
+ 751.000001n V_hig
+ 751.100000n V_hig
+ 751.100001n V_hig
+ 751.200000n V_hig
+ 751.200001n V_hig
+ 751.300000n V_hig
+ 751.300001n V_hig
+ 751.400000n V_hig
+ 751.400001n V_hig
+ 751.500000n V_hig
+ 751.500001n V_hig
+ 751.600000n V_hig
+ 751.600001n V_hig
+ 751.700000n V_hig
+ 751.700001n V_hig
+ 751.800000n V_hig
+ 751.800001n V_hig
+ 751.900000n V_hig
+ 751.900001n V_hig
+ 752.000000n V_hig
+ 752.000001n V_low
+ 752.100000n V_low
+ 752.100001n V_low
+ 752.200000n V_low
+ 752.200001n V_low
+ 752.300000n V_low
+ 752.300001n V_low
+ 752.400000n V_low
+ 752.400001n V_low
+ 752.500000n V_low
+ 752.500001n V_low
+ 752.600000n V_low
+ 752.600001n V_low
+ 752.700000n V_low
+ 752.700001n V_low
+ 752.800000n V_low
+ 752.800001n V_low
+ 752.900000n V_low
+ 752.900001n V_low
+ 753.000000n V_low
+ 753.000001n V_hig
+ 753.100000n V_hig
+ 753.100001n V_hig
+ 753.200000n V_hig
+ 753.200001n V_hig
+ 753.300000n V_hig
+ 753.300001n V_hig
+ 753.400000n V_hig
+ 753.400001n V_hig
+ 753.500000n V_hig
+ 753.500001n V_hig
+ 753.600000n V_hig
+ 753.600001n V_hig
+ 753.700000n V_hig
+ 753.700001n V_hig
+ 753.800000n V_hig
+ 753.800001n V_hig
+ 753.900000n V_hig
+ 753.900001n V_hig
+ 754.000000n V_hig
+ 754.000001n V_low
+ 754.100000n V_low
+ 754.100001n V_low
+ 754.200000n V_low
+ 754.200001n V_low
+ 754.300000n V_low
+ 754.300001n V_low
+ 754.400000n V_low
+ 754.400001n V_low
+ 754.500000n V_low
+ 754.500001n V_low
+ 754.600000n V_low
+ 754.600001n V_low
+ 754.700000n V_low
+ 754.700001n V_low
+ 754.800000n V_low
+ 754.800001n V_low
+ 754.900000n V_low
+ 754.900001n V_low
+ 755.000000n V_low
+ 755.000001n V_hig
+ 755.100000n V_hig
+ 755.100001n V_hig
+ 755.200000n V_hig
+ 755.200001n V_hig
+ 755.300000n V_hig
+ 755.300001n V_hig
+ 755.400000n V_hig
+ 755.400001n V_hig
+ 755.500000n V_hig
+ 755.500001n V_hig
+ 755.600000n V_hig
+ 755.600001n V_hig
+ 755.700000n V_hig
+ 755.700001n V_hig
+ 755.800000n V_hig
+ 755.800001n V_hig
+ 755.900000n V_hig
+ 755.900001n V_hig
+ 756.000000n V_hig
+ 756.000001n V_low
+ 756.100000n V_low
+ 756.100001n V_low
+ 756.200000n V_low
+ 756.200001n V_low
+ 756.300000n V_low
+ 756.300001n V_low
+ 756.400000n V_low
+ 756.400001n V_low
+ 756.500000n V_low
+ 756.500001n V_low
+ 756.600000n V_low
+ 756.600001n V_low
+ 756.700000n V_low
+ 756.700001n V_low
+ 756.800000n V_low
+ 756.800001n V_low
+ 756.900000n V_low
+ 756.900001n V_low
+ 757.000000n V_low
+ 757.000001n V_low
+ 757.100000n V_low
+ 757.100001n V_low
+ 757.200000n V_low
+ 757.200001n V_low
+ 757.300000n V_low
+ 757.300001n V_low
+ 757.400000n V_low
+ 757.400001n V_low
+ 757.500000n V_low
+ 757.500001n V_low
+ 757.600000n V_low
+ 757.600001n V_low
+ 757.700000n V_low
+ 757.700001n V_low
+ 757.800000n V_low
+ 757.800001n V_low
+ 757.900000n V_low
+ 757.900001n V_low
+ 758.000000n V_low
+ 758.000001n V_low
+ 758.100000n V_low
+ 758.100001n V_low
+ 758.200000n V_low
+ 758.200001n V_low
+ 758.300000n V_low
+ 758.300001n V_low
+ 758.400000n V_low
+ 758.400001n V_low
+ 758.500000n V_low
+ 758.500001n V_low
+ 758.600000n V_low
+ 758.600001n V_low
+ 758.700000n V_low
+ 758.700001n V_low
+ 758.800000n V_low
+ 758.800001n V_low
+ 758.900000n V_low
+ 758.900001n V_low
+ 759.000000n V_low
+ 759.000001n V_hig
+ 759.100000n V_hig
+ 759.100001n V_hig
+ 759.200000n V_hig
+ 759.200001n V_hig
+ 759.300000n V_hig
+ 759.300001n V_hig
+ 759.400000n V_hig
+ 759.400001n V_hig
+ 759.500000n V_hig
+ 759.500001n V_hig
+ 759.600000n V_hig
+ 759.600001n V_hig
+ 759.700000n V_hig
+ 759.700001n V_hig
+ 759.800000n V_hig
+ 759.800001n V_hig
+ 759.900000n V_hig
+ 759.900001n V_hig
+ 760.000000n V_hig
+ 760.000001n V_low
+ 760.100000n V_low
+ 760.100001n V_low
+ 760.200000n V_low
+ 760.200001n V_low
+ 760.300000n V_low
+ 760.300001n V_low
+ 760.400000n V_low
+ 760.400001n V_low
+ 760.500000n V_low
+ 760.500001n V_low
+ 760.600000n V_low
+ 760.600001n V_low
+ 760.700000n V_low
+ 760.700001n V_low
+ 760.800000n V_low
+ 760.800001n V_low
+ 760.900000n V_low
+ 760.900001n V_low
+ 761.000000n V_low
+ 761.000001n V_hig
+ 761.100000n V_hig
+ 761.100001n V_hig
+ 761.200000n V_hig
+ 761.200001n V_hig
+ 761.300000n V_hig
+ 761.300001n V_hig
+ 761.400000n V_hig
+ 761.400001n V_hig
+ 761.500000n V_hig
+ 761.500001n V_hig
+ 761.600000n V_hig
+ 761.600001n V_hig
+ 761.700000n V_hig
+ 761.700001n V_hig
+ 761.800000n V_hig
+ 761.800001n V_hig
+ 761.900000n V_hig
+ 761.900001n V_hig
+ 762.000000n V_hig
+ 762.000001n V_low
+ 762.100000n V_low
+ 762.100001n V_low
+ 762.200000n V_low
+ 762.200001n V_low
+ 762.300000n V_low
+ 762.300001n V_low
+ 762.400000n V_low
+ 762.400001n V_low
+ 762.500000n V_low
+ 762.500001n V_low
+ 762.600000n V_low
+ 762.600001n V_low
+ 762.700000n V_low
+ 762.700001n V_low
+ 762.800000n V_low
+ 762.800001n V_low
+ 762.900000n V_low
+ 762.900001n V_low
+ 763.000000n V_low
+ 763.000001n V_hig
+ 763.100000n V_hig
+ 763.100001n V_hig
+ 763.200000n V_hig
+ 763.200001n V_hig
+ 763.300000n V_hig
+ 763.300001n V_hig
+ 763.400000n V_hig
+ 763.400001n V_hig
+ 763.500000n V_hig
+ 763.500001n V_hig
+ 763.600000n V_hig
+ 763.600001n V_hig
+ 763.700000n V_hig
+ 763.700001n V_hig
+ 763.800000n V_hig
+ 763.800001n V_hig
+ 763.900000n V_hig
+ 763.900001n V_hig
+ 764.000000n V_hig
+ 764.000001n V_low
+ 764.100000n V_low
+ 764.100001n V_low
+ 764.200000n V_low
+ 764.200001n V_low
+ 764.300000n V_low
+ 764.300001n V_low
+ 764.400000n V_low
+ 764.400001n V_low
+ 764.500000n V_low
+ 764.500001n V_low
+ 764.600000n V_low
+ 764.600001n V_low
+ 764.700000n V_low
+ 764.700001n V_low
+ 764.800000n V_low
+ 764.800001n V_low
+ 764.900000n V_low
+ 764.900001n V_low
+ 765.000000n V_low
+ 765.000001n V_low
+ 765.100000n V_low
+ 765.100001n V_low
+ 765.200000n V_low
+ 765.200001n V_low
+ 765.300000n V_low
+ 765.300001n V_low
+ 765.400000n V_low
+ 765.400001n V_low
+ 765.500000n V_low
+ 765.500001n V_low
+ 765.600000n V_low
+ 765.600001n V_low
+ 765.700000n V_low
+ 765.700001n V_low
+ 765.800000n V_low
+ 765.800001n V_low
+ 765.900000n V_low
+ 765.900001n V_low
+ 766.000000n V_low
+ 766.000001n V_low
+ 766.100000n V_low
+ 766.100001n V_low
+ 766.200000n V_low
+ 766.200001n V_low
+ 766.300000n V_low
+ 766.300001n V_low
+ 766.400000n V_low
+ 766.400001n V_low
+ 766.500000n V_low
+ 766.500001n V_low
+ 766.600000n V_low
+ 766.600001n V_low
+ 766.700000n V_low
+ 766.700001n V_low
+ 766.800000n V_low
+ 766.800001n V_low
+ 766.900000n V_low
+ 766.900001n V_low
+ 767.000000n V_low
+ 767.000001n V_hig
+ 767.100000n V_hig
+ 767.100001n V_hig
+ 767.200000n V_hig
+ 767.200001n V_hig
+ 767.300000n V_hig
+ 767.300001n V_hig
+ 767.400000n V_hig
+ 767.400001n V_hig
+ 767.500000n V_hig
+ 767.500001n V_hig
+ 767.600000n V_hig
+ 767.600001n V_hig
+ 767.700000n V_hig
+ 767.700001n V_hig
+ 767.800000n V_hig
+ 767.800001n V_hig
+ 767.900000n V_hig
+ 767.900001n V_hig
+ 768.000000n V_hig
+ 768.000001n V_low
+ 768.100000n V_low
+ 768.100001n V_low
+ 768.200000n V_low
+ 768.200001n V_low
+ 768.300000n V_low
+ 768.300001n V_low
+ 768.400000n V_low
+ 768.400001n V_low
+ 768.500000n V_low
+ 768.500001n V_low
+ 768.600000n V_low
+ 768.600001n V_low
+ 768.700000n V_low
+ 768.700001n V_low
+ 768.800000n V_low
+ 768.800001n V_low
+ 768.900000n V_low
+ 768.900001n V_low
+ 769.000000n V_low
+ 769.000001n V_hig
+ 769.100000n V_hig
+ 769.100001n V_hig
+ 769.200000n V_hig
+ 769.200001n V_hig
+ 769.300000n V_hig
+ 769.300001n V_hig
+ 769.400000n V_hig
+ 769.400001n V_hig
+ 769.500000n V_hig
+ 769.500001n V_hig
+ 769.600000n V_hig
+ 769.600001n V_hig
+ 769.700000n V_hig
+ 769.700001n V_hig
+ 769.800000n V_hig
+ 769.800001n V_hig
+ 769.900000n V_hig
+ 769.900001n V_hig
+ 770.000000n V_hig
+ 770.000001n V_hig
+ 770.100000n V_hig
+ 770.100001n V_hig
+ 770.200000n V_hig
+ 770.200001n V_hig
+ 770.300000n V_hig
+ 770.300001n V_hig
+ 770.400000n V_hig
+ 770.400001n V_hig
+ 770.500000n V_hig
+ 770.500001n V_hig
+ 770.600000n V_hig
+ 770.600001n V_hig
+ 770.700000n V_hig
+ 770.700001n V_hig
+ 770.800000n V_hig
+ 770.800001n V_hig
+ 770.900000n V_hig
+ 770.900001n V_hig
+ 771.000000n V_hig
+ 771.000001n V_low
+ 771.100000n V_low
+ 771.100001n V_low
+ 771.200000n V_low
+ 771.200001n V_low
+ 771.300000n V_low
+ 771.300001n V_low
+ 771.400000n V_low
+ 771.400001n V_low
+ 771.500000n V_low
+ 771.500001n V_low
+ 771.600000n V_low
+ 771.600001n V_low
+ 771.700000n V_low
+ 771.700001n V_low
+ 771.800000n V_low
+ 771.800001n V_low
+ 771.900000n V_low
+ 771.900001n V_low
+ 772.000000n V_low
+ 772.000001n V_hig
+ 772.100000n V_hig
+ 772.100001n V_hig
+ 772.200000n V_hig
+ 772.200001n V_hig
+ 772.300000n V_hig
+ 772.300001n V_hig
+ 772.400000n V_hig
+ 772.400001n V_hig
+ 772.500000n V_hig
+ 772.500001n V_hig
+ 772.600000n V_hig
+ 772.600001n V_hig
+ 772.700000n V_hig
+ 772.700001n V_hig
+ 772.800000n V_hig
+ 772.800001n V_hig
+ 772.900000n V_hig
+ 772.900001n V_hig
+ 773.000000n V_hig
+ 773.000001n V_low
+ 773.100000n V_low
+ 773.100001n V_low
+ 773.200000n V_low
+ 773.200001n V_low
+ 773.300000n V_low
+ 773.300001n V_low
+ 773.400000n V_low
+ 773.400001n V_low
+ 773.500000n V_low
+ 773.500001n V_low
+ 773.600000n V_low
+ 773.600001n V_low
+ 773.700000n V_low
+ 773.700001n V_low
+ 773.800000n V_low
+ 773.800001n V_low
+ 773.900000n V_low
+ 773.900001n V_low
+ 774.000000n V_low
+ 774.000001n V_hig
+ 774.100000n V_hig
+ 774.100001n V_hig
+ 774.200000n V_hig
+ 774.200001n V_hig
+ 774.300000n V_hig
+ 774.300001n V_hig
+ 774.400000n V_hig
+ 774.400001n V_hig
+ 774.500000n V_hig
+ 774.500001n V_hig
+ 774.600000n V_hig
+ 774.600001n V_hig
+ 774.700000n V_hig
+ 774.700001n V_hig
+ 774.800000n V_hig
+ 774.800001n V_hig
+ 774.900000n V_hig
+ 774.900001n V_hig
+ 775.000000n V_hig
+ 775.000001n V_low
+ 775.100000n V_low
+ 775.100001n V_low
+ 775.200000n V_low
+ 775.200001n V_low
+ 775.300000n V_low
+ 775.300001n V_low
+ 775.400000n V_low
+ 775.400001n V_low
+ 775.500000n V_low
+ 775.500001n V_low
+ 775.600000n V_low
+ 775.600001n V_low
+ 775.700000n V_low
+ 775.700001n V_low
+ 775.800000n V_low
+ 775.800001n V_low
+ 775.900000n V_low
+ 775.900001n V_low
+ 776.000000n V_low
+ 776.000001n V_hig
+ 776.100000n V_hig
+ 776.100001n V_hig
+ 776.200000n V_hig
+ 776.200001n V_hig
+ 776.300000n V_hig
+ 776.300001n V_hig
+ 776.400000n V_hig
+ 776.400001n V_hig
+ 776.500000n V_hig
+ 776.500001n V_hig
+ 776.600000n V_hig
+ 776.600001n V_hig
+ 776.700000n V_hig
+ 776.700001n V_hig
+ 776.800000n V_hig
+ 776.800001n V_hig
+ 776.900000n V_hig
+ 776.900001n V_hig
+ 777.000000n V_hig
+ 777.000001n V_low
+ 777.100000n V_low
+ 777.100001n V_low
+ 777.200000n V_low
+ 777.200001n V_low
+ 777.300000n V_low
+ 777.300001n V_low
+ 777.400000n V_low
+ 777.400001n V_low
+ 777.500000n V_low
+ 777.500001n V_low
+ 777.600000n V_low
+ 777.600001n V_low
+ 777.700000n V_low
+ 777.700001n V_low
+ 777.800000n V_low
+ 777.800001n V_low
+ 777.900000n V_low
+ 777.900001n V_low
+ 778.000000n V_low
+ 778.000001n V_hig
+ 778.100000n V_hig
+ 778.100001n V_hig
+ 778.200000n V_hig
+ 778.200001n V_hig
+ 778.300000n V_hig
+ 778.300001n V_hig
+ 778.400000n V_hig
+ 778.400001n V_hig
+ 778.500000n V_hig
+ 778.500001n V_hig
+ 778.600000n V_hig
+ 778.600001n V_hig
+ 778.700000n V_hig
+ 778.700001n V_hig
+ 778.800000n V_hig
+ 778.800001n V_hig
+ 778.900000n V_hig
+ 778.900001n V_hig
+ 779.000000n V_hig
+ 779.000001n V_hig
+ 779.100000n V_hig
+ 779.100001n V_hig
+ 779.200000n V_hig
+ 779.200001n V_hig
+ 779.300000n V_hig
+ 779.300001n V_hig
+ 779.400000n V_hig
+ 779.400001n V_hig
+ 779.500000n V_hig
+ 779.500001n V_hig
+ 779.600000n V_hig
+ 779.600001n V_hig
+ 779.700000n V_hig
+ 779.700001n V_hig
+ 779.800000n V_hig
+ 779.800001n V_hig
+ 779.900000n V_hig
+ 779.900001n V_hig
+ 780.000000n V_hig
+ 780.000001n V_low
+ 780.100000n V_low
+ 780.100001n V_low
+ 780.200000n V_low
+ 780.200001n V_low
+ 780.300000n V_low
+ 780.300001n V_low
+ 780.400000n V_low
+ 780.400001n V_low
+ 780.500000n V_low
+ 780.500001n V_low
+ 780.600000n V_low
+ 780.600001n V_low
+ 780.700000n V_low
+ 780.700001n V_low
+ 780.800000n V_low
+ 780.800001n V_low
+ 780.900000n V_low
+ 780.900001n V_low
+ 781.000000n V_low
+ 781.000001n V_hig
+ 781.100000n V_hig
+ 781.100001n V_hig
+ 781.200000n V_hig
+ 781.200001n V_hig
+ 781.300000n V_hig
+ 781.300001n V_hig
+ 781.400000n V_hig
+ 781.400001n V_hig
+ 781.500000n V_hig
+ 781.500001n V_hig
+ 781.600000n V_hig
+ 781.600001n V_hig
+ 781.700000n V_hig
+ 781.700001n V_hig
+ 781.800000n V_hig
+ 781.800001n V_hig
+ 781.900000n V_hig
+ 781.900001n V_hig
+ 782.000000n V_hig
+ 782.000001n V_hig
+ 782.100000n V_hig
+ 782.100001n V_hig
+ 782.200000n V_hig
+ 782.200001n V_hig
+ 782.300000n V_hig
+ 782.300001n V_hig
+ 782.400000n V_hig
+ 782.400001n V_hig
+ 782.500000n V_hig
+ 782.500001n V_hig
+ 782.600000n V_hig
+ 782.600001n V_hig
+ 782.700000n V_hig
+ 782.700001n V_hig
+ 782.800000n V_hig
+ 782.800001n V_hig
+ 782.900000n V_hig
+ 782.900001n V_hig
+ 783.000000n V_hig
+ 783.000001n V_hig
+ 783.100000n V_hig
+ 783.100001n V_hig
+ 783.200000n V_hig
+ 783.200001n V_hig
+ 783.300000n V_hig
+ 783.300001n V_hig
+ 783.400000n V_hig
+ 783.400001n V_hig
+ 783.500000n V_hig
+ 783.500001n V_hig
+ 783.600000n V_hig
+ 783.600001n V_hig
+ 783.700000n V_hig
+ 783.700001n V_hig
+ 783.800000n V_hig
+ 783.800001n V_hig
+ 783.900000n V_hig
+ 783.900001n V_hig
+ 784.000000n V_hig
+ 784.000001n V_low
+ 784.100000n V_low
+ 784.100001n V_low
+ 784.200000n V_low
+ 784.200001n V_low
+ 784.300000n V_low
+ 784.300001n V_low
+ 784.400000n V_low
+ 784.400001n V_low
+ 784.500000n V_low
+ 784.500001n V_low
+ 784.600000n V_low
+ 784.600001n V_low
+ 784.700000n V_low
+ 784.700001n V_low
+ 784.800000n V_low
+ 784.800001n V_low
+ 784.900000n V_low
+ 784.900001n V_low
+ 785.000000n V_low
+ 785.000001n V_hig
+ 785.100000n V_hig
+ 785.100001n V_hig
+ 785.200000n V_hig
+ 785.200001n V_hig
+ 785.300000n V_hig
+ 785.300001n V_hig
+ 785.400000n V_hig
+ 785.400001n V_hig
+ 785.500000n V_hig
+ 785.500001n V_hig
+ 785.600000n V_hig
+ 785.600001n V_hig
+ 785.700000n V_hig
+ 785.700001n V_hig
+ 785.800000n V_hig
+ 785.800001n V_hig
+ 785.900000n V_hig
+ 785.900001n V_hig
+ 786.000000n V_hig
+ 786.000001n V_low
+ 786.100000n V_low
+ 786.100001n V_low
+ 786.200000n V_low
+ 786.200001n V_low
+ 786.300000n V_low
+ 786.300001n V_low
+ 786.400000n V_low
+ 786.400001n V_low
+ 786.500000n V_low
+ 786.500001n V_low
+ 786.600000n V_low
+ 786.600001n V_low
+ 786.700000n V_low
+ 786.700001n V_low
+ 786.800000n V_low
+ 786.800001n V_low
+ 786.900000n V_low
+ 786.900001n V_low
+ 787.000000n V_low
+ 787.000001n V_low
+ 787.100000n V_low
+ 787.100001n V_low
+ 787.200000n V_low
+ 787.200001n V_low
+ 787.300000n V_low
+ 787.300001n V_low
+ 787.400000n V_low
+ 787.400001n V_low
+ 787.500000n V_low
+ 787.500001n V_low
+ 787.600000n V_low
+ 787.600001n V_low
+ 787.700000n V_low
+ 787.700001n V_low
+ 787.800000n V_low
+ 787.800001n V_low
+ 787.900000n V_low
+ 787.900001n V_low
+ 788.000000n V_low
+ 788.000001n V_low
+ 788.100000n V_low
+ 788.100001n V_low
+ 788.200000n V_low
+ 788.200001n V_low
+ 788.300000n V_low
+ 788.300001n V_low
+ 788.400000n V_low
+ 788.400001n V_low
+ 788.500000n V_low
+ 788.500001n V_low
+ 788.600000n V_low
+ 788.600001n V_low
+ 788.700000n V_low
+ 788.700001n V_low
+ 788.800000n V_low
+ 788.800001n V_low
+ 788.900000n V_low
+ 788.900001n V_low
+ 789.000000n V_low
+ 789.000001n V_low
+ 789.100000n V_low
+ 789.100001n V_low
+ 789.200000n V_low
+ 789.200001n V_low
+ 789.300000n V_low
+ 789.300001n V_low
+ 789.400000n V_low
+ 789.400001n V_low
+ 789.500000n V_low
+ 789.500001n V_low
+ 789.600000n V_low
+ 789.600001n V_low
+ 789.700000n V_low
+ 789.700001n V_low
+ 789.800000n V_low
+ 789.800001n V_low
+ 789.900000n V_low
+ 789.900001n V_low
+ 790.000000n V_low
+ 790.000001n V_hig
+ 790.100000n V_hig
+ 790.100001n V_hig
+ 790.200000n V_hig
+ 790.200001n V_hig
+ 790.300000n V_hig
+ 790.300001n V_hig
+ 790.400000n V_hig
+ 790.400001n V_hig
+ 790.500000n V_hig
+ 790.500001n V_hig
+ 790.600000n V_hig
+ 790.600001n V_hig
+ 790.700000n V_hig
+ 790.700001n V_hig
+ 790.800000n V_hig
+ 790.800001n V_hig
+ 790.900000n V_hig
+ 790.900001n V_hig
+ 791.000000n V_hig
+ 791.000001n V_low
+ 791.100000n V_low
+ 791.100001n V_low
+ 791.200000n V_low
+ 791.200001n V_low
+ 791.300000n V_low
+ 791.300001n V_low
+ 791.400000n V_low
+ 791.400001n V_low
+ 791.500000n V_low
+ 791.500001n V_low
+ 791.600000n V_low
+ 791.600001n V_low
+ 791.700000n V_low
+ 791.700001n V_low
+ 791.800000n V_low
+ 791.800001n V_low
+ 791.900000n V_low
+ 791.900001n V_low
+ 792.000000n V_low
+ 792.000001n V_hig
+ 792.100000n V_hig
+ 792.100001n V_hig
+ 792.200000n V_hig
+ 792.200001n V_hig
+ 792.300000n V_hig
+ 792.300001n V_hig
+ 792.400000n V_hig
+ 792.400001n V_hig
+ 792.500000n V_hig
+ 792.500001n V_hig
+ 792.600000n V_hig
+ 792.600001n V_hig
+ 792.700000n V_hig
+ 792.700001n V_hig
+ 792.800000n V_hig
+ 792.800001n V_hig
+ 792.900000n V_hig
+ 792.900001n V_hig
+ 793.000000n V_hig
+ 793.000001n V_hig
+ 793.100000n V_hig
+ 793.100001n V_hig
+ 793.200000n V_hig
+ 793.200001n V_hig
+ 793.300000n V_hig
+ 793.300001n V_hig
+ 793.400000n V_hig
+ 793.400001n V_hig
+ 793.500000n V_hig
+ 793.500001n V_hig
+ 793.600000n V_hig
+ 793.600001n V_hig
+ 793.700000n V_hig
+ 793.700001n V_hig
+ 793.800000n V_hig
+ 793.800001n V_hig
+ 793.900000n V_hig
+ 793.900001n V_hig
+ 794.000000n V_hig
+ 794.000001n V_low
+ 794.100000n V_low
+ 794.100001n V_low
+ 794.200000n V_low
+ 794.200001n V_low
+ 794.300000n V_low
+ 794.300001n V_low
+ 794.400000n V_low
+ 794.400001n V_low
+ 794.500000n V_low
+ 794.500001n V_low
+ 794.600000n V_low
+ 794.600001n V_low
+ 794.700000n V_low
+ 794.700001n V_low
+ 794.800000n V_low
+ 794.800001n V_low
+ 794.900000n V_low
+ 794.900001n V_low
+ 795.000000n V_low
+ 795.000001n V_hig
+ 795.100000n V_hig
+ 795.100001n V_hig
+ 795.200000n V_hig
+ 795.200001n V_hig
+ 795.300000n V_hig
+ 795.300001n V_hig
+ 795.400000n V_hig
+ 795.400001n V_hig
+ 795.500000n V_hig
+ 795.500001n V_hig
+ 795.600000n V_hig
+ 795.600001n V_hig
+ 795.700000n V_hig
+ 795.700001n V_hig
+ 795.800000n V_hig
+ 795.800001n V_hig
+ 795.900000n V_hig
+ 795.900001n V_hig
+ 796.000000n V_hig
+ 796.000001n V_low
+ 796.100000n V_low
+ 796.100001n V_low
+ 796.200000n V_low
+ 796.200001n V_low
+ 796.300000n V_low
+ 796.300001n V_low
+ 796.400000n V_low
+ 796.400001n V_low
+ 796.500000n V_low
+ 796.500001n V_low
+ 796.600000n V_low
+ 796.600001n V_low
+ 796.700000n V_low
+ 796.700001n V_low
+ 796.800000n V_low
+ 796.800001n V_low
+ 796.900000n V_low
+ 796.900001n V_low
+ 797.000000n V_low
+ 797.000001n V_hig
+ 797.100000n V_hig
+ 797.100001n V_hig
+ 797.200000n V_hig
+ 797.200001n V_hig
+ 797.300000n V_hig
+ 797.300001n V_hig
+ 797.400000n V_hig
+ 797.400001n V_hig
+ 797.500000n V_hig
+ 797.500001n V_hig
+ 797.600000n V_hig
+ 797.600001n V_hig
+ 797.700000n V_hig
+ 797.700001n V_hig
+ 797.800000n V_hig
+ 797.800001n V_hig
+ 797.900000n V_hig
+ 797.900001n V_hig
+ 798.000000n V_hig
+ 798.000001n V_low
+ 798.100000n V_low
+ 798.100001n V_low
+ 798.200000n V_low
+ 798.200001n V_low
+ 798.300000n V_low
+ 798.300001n V_low
+ 798.400000n V_low
+ 798.400001n V_low
+ 798.500000n V_low
+ 798.500001n V_low
+ 798.600000n V_low
+ 798.600001n V_low
+ 798.700000n V_low
+ 798.700001n V_low
+ 798.800000n V_low
+ 798.800001n V_low
+ 798.900000n V_low
+ 798.900001n V_low
+ 799.000000n V_low
+ 799.000001n V_low
+ 799.100000n V_low
+ 799.100001n V_low
+ 799.200000n V_low
+ 799.200001n V_low
+ 799.300000n V_low
+ 799.300001n V_low
+ 799.400000n V_low
+ 799.400001n V_low
+ 799.500000n V_low
+ 799.500001n V_low
+ 799.600000n V_low
+ 799.600001n V_low
+ 799.700000n V_low
+ 799.700001n V_low
+ 799.800000n V_low
+ 799.800001n V_low
+ 799.900000n V_low
+ 799.900001n V_low
+ 800.000000n V_low
+ 800.000001n V_low
+ 800.100000n V_low
+ 800.100001n V_low
+ 800.200000n V_low
+ 800.200001n V_low
+ 800.300000n V_low
+ 800.300001n V_low
+ 800.400000n V_low
+ 800.400001n V_low
+ 800.500000n V_low
+ 800.500001n V_low
+ 800.600000n V_low
+ 800.600001n V_low
+ 800.700000n V_low
+ 800.700001n V_low
+ 800.800000n V_low
+ 800.800001n V_low
+ 800.900000n V_low
+ 800.900001n V_low
+ 801.000000n V_low
+ 801.000001n V_hig
+ 801.100000n V_hig
+ 801.100001n V_hig
+ 801.200000n V_hig
+ 801.200001n V_hig
+ 801.300000n V_hig
+ 801.300001n V_hig
+ 801.400000n V_hig
+ 801.400001n V_hig
+ 801.500000n V_hig
+ 801.500001n V_hig
+ 801.600000n V_hig
+ 801.600001n V_hig
+ 801.700000n V_hig
+ 801.700001n V_hig
+ 801.800000n V_hig
+ 801.800001n V_hig
+ 801.900000n V_hig
+ 801.900001n V_hig
+ 802.000000n V_hig
+ 802.000001n V_low
+ 802.100000n V_low
+ 802.100001n V_low
+ 802.200000n V_low
+ 802.200001n V_low
+ 802.300000n V_low
+ 802.300001n V_low
+ 802.400000n V_low
+ 802.400001n V_low
+ 802.500000n V_low
+ 802.500001n V_low
+ 802.600000n V_low
+ 802.600001n V_low
+ 802.700000n V_low
+ 802.700001n V_low
+ 802.800000n V_low
+ 802.800001n V_low
+ 802.900000n V_low
+ 802.900001n V_low
+ 803.000000n V_low
+ 803.000001n V_low
+ 803.100000n V_low
+ 803.100001n V_low
+ 803.200000n V_low
+ 803.200001n V_low
+ 803.300000n V_low
+ 803.300001n V_low
+ 803.400000n V_low
+ 803.400001n V_low
+ 803.500000n V_low
+ 803.500001n V_low
+ 803.600000n V_low
+ 803.600001n V_low
+ 803.700000n V_low
+ 803.700001n V_low
+ 803.800000n V_low
+ 803.800001n V_low
+ 803.900000n V_low
+ 803.900001n V_low
+ 804.000000n V_low
+ 804.000001n V_low
+ 804.100000n V_low
+ 804.100001n V_low
+ 804.200000n V_low
+ 804.200001n V_low
+ 804.300000n V_low
+ 804.300001n V_low
+ 804.400000n V_low
+ 804.400001n V_low
+ 804.500000n V_low
+ 804.500001n V_low
+ 804.600000n V_low
+ 804.600001n V_low
+ 804.700000n V_low
+ 804.700001n V_low
+ 804.800000n V_low
+ 804.800001n V_low
+ 804.900000n V_low
+ 804.900001n V_low
+ 805.000000n V_low
+ 805.000001n V_hig
+ 805.100000n V_hig
+ 805.100001n V_hig
+ 805.200000n V_hig
+ 805.200001n V_hig
+ 805.300000n V_hig
+ 805.300001n V_hig
+ 805.400000n V_hig
+ 805.400001n V_hig
+ 805.500000n V_hig
+ 805.500001n V_hig
+ 805.600000n V_hig
+ 805.600001n V_hig
+ 805.700000n V_hig
+ 805.700001n V_hig
+ 805.800000n V_hig
+ 805.800001n V_hig
+ 805.900000n V_hig
+ 805.900001n V_hig
+ 806.000000n V_hig
+ 806.000001n V_hig
+ 806.100000n V_hig
+ 806.100001n V_hig
+ 806.200000n V_hig
+ 806.200001n V_hig
+ 806.300000n V_hig
+ 806.300001n V_hig
+ 806.400000n V_hig
+ 806.400001n V_hig
+ 806.500000n V_hig
+ 806.500001n V_hig
+ 806.600000n V_hig
+ 806.600001n V_hig
+ 806.700000n V_hig
+ 806.700001n V_hig
+ 806.800000n V_hig
+ 806.800001n V_hig
+ 806.900000n V_hig
+ 806.900001n V_hig
+ 807.000000n V_hig
+ 807.000001n V_low
+ 807.100000n V_low
+ 807.100001n V_low
+ 807.200000n V_low
+ 807.200001n V_low
+ 807.300000n V_low
+ 807.300001n V_low
+ 807.400000n V_low
+ 807.400001n V_low
+ 807.500000n V_low
+ 807.500001n V_low
+ 807.600000n V_low
+ 807.600001n V_low
+ 807.700000n V_low
+ 807.700001n V_low
+ 807.800000n V_low
+ 807.800001n V_low
+ 807.900000n V_low
+ 807.900001n V_low
+ 808.000000n V_low
+ 808.000001n V_low
+ 808.100000n V_low
+ 808.100001n V_low
+ 808.200000n V_low
+ 808.200001n V_low
+ 808.300000n V_low
+ 808.300001n V_low
+ 808.400000n V_low
+ 808.400001n V_low
+ 808.500000n V_low
+ 808.500001n V_low
+ 808.600000n V_low
+ 808.600001n V_low
+ 808.700000n V_low
+ 808.700001n V_low
+ 808.800000n V_low
+ 808.800001n V_low
+ 808.900000n V_low
+ 808.900001n V_low
+ 809.000000n V_low
+ 809.000001n V_low
+ 809.100000n V_low
+ 809.100001n V_low
+ 809.200000n V_low
+ 809.200001n V_low
+ 809.300000n V_low
+ 809.300001n V_low
+ 809.400000n V_low
+ 809.400001n V_low
+ 809.500000n V_low
+ 809.500001n V_low
+ 809.600000n V_low
+ 809.600001n V_low
+ 809.700000n V_low
+ 809.700001n V_low
+ 809.800000n V_low
+ 809.800001n V_low
+ 809.900000n V_low
+ 809.900001n V_low
+ 810.000000n V_low
+ 810.000001n V_low
+ 810.100000n V_low
+ 810.100001n V_low
+ 810.200000n V_low
+ 810.200001n V_low
+ 810.300000n V_low
+ 810.300001n V_low
+ 810.400000n V_low
+ 810.400001n V_low
+ 810.500000n V_low
+ 810.500001n V_low
+ 810.600000n V_low
+ 810.600001n V_low
+ 810.700000n V_low
+ 810.700001n V_low
+ 810.800000n V_low
+ 810.800001n V_low
+ 810.900000n V_low
+ 810.900001n V_low
+ 811.000000n V_low
+ 811.000001n V_low
+ 811.100000n V_low
+ 811.100001n V_low
+ 811.200000n V_low
+ 811.200001n V_low
+ 811.300000n V_low
+ 811.300001n V_low
+ 811.400000n V_low
+ 811.400001n V_low
+ 811.500000n V_low
+ 811.500001n V_low
+ 811.600000n V_low
+ 811.600001n V_low
+ 811.700000n V_low
+ 811.700001n V_low
+ 811.800000n V_low
+ 811.800001n V_low
+ 811.900000n V_low
+ 811.900001n V_low
+ 812.000000n V_low
+ 812.000001n V_low
+ 812.100000n V_low
+ 812.100001n V_low
+ 812.200000n V_low
+ 812.200001n V_low
+ 812.300000n V_low
+ 812.300001n V_low
+ 812.400000n V_low
+ 812.400001n V_low
+ 812.500000n V_low
+ 812.500001n V_low
+ 812.600000n V_low
+ 812.600001n V_low
+ 812.700000n V_low
+ 812.700001n V_low
+ 812.800000n V_low
+ 812.800001n V_low
+ 812.900000n V_low
+ 812.900001n V_low
+ 813.000000n V_low
+ 813.000001n V_hig
+ 813.100000n V_hig
+ 813.100001n V_hig
+ 813.200000n V_hig
+ 813.200001n V_hig
+ 813.300000n V_hig
+ 813.300001n V_hig
+ 813.400000n V_hig
+ 813.400001n V_hig
+ 813.500000n V_hig
+ 813.500001n V_hig
+ 813.600000n V_hig
+ 813.600001n V_hig
+ 813.700000n V_hig
+ 813.700001n V_hig
+ 813.800000n V_hig
+ 813.800001n V_hig
+ 813.900000n V_hig
+ 813.900001n V_hig
+ 814.000000n V_hig
+ 814.000001n V_low
+ 814.100000n V_low
+ 814.100001n V_low
+ 814.200000n V_low
+ 814.200001n V_low
+ 814.300000n V_low
+ 814.300001n V_low
+ 814.400000n V_low
+ 814.400001n V_low
+ 814.500000n V_low
+ 814.500001n V_low
+ 814.600000n V_low
+ 814.600001n V_low
+ 814.700000n V_low
+ 814.700001n V_low
+ 814.800000n V_low
+ 814.800001n V_low
+ 814.900000n V_low
+ 814.900001n V_low
+ 815.000000n V_low
+ 815.000001n V_hig
+ 815.100000n V_hig
+ 815.100001n V_hig
+ 815.200000n V_hig
+ 815.200001n V_hig
+ 815.300000n V_hig
+ 815.300001n V_hig
+ 815.400000n V_hig
+ 815.400001n V_hig
+ 815.500000n V_hig
+ 815.500001n V_hig
+ 815.600000n V_hig
+ 815.600001n V_hig
+ 815.700000n V_hig
+ 815.700001n V_hig
+ 815.800000n V_hig
+ 815.800001n V_hig
+ 815.900000n V_hig
+ 815.900001n V_hig
+ 816.000000n V_hig
+ 816.000001n V_low
+ 816.100000n V_low
+ 816.100001n V_low
+ 816.200000n V_low
+ 816.200001n V_low
+ 816.300000n V_low
+ 816.300001n V_low
+ 816.400000n V_low
+ 816.400001n V_low
+ 816.500000n V_low
+ 816.500001n V_low
+ 816.600000n V_low
+ 816.600001n V_low
+ 816.700000n V_low
+ 816.700001n V_low
+ 816.800000n V_low
+ 816.800001n V_low
+ 816.900000n V_low
+ 816.900001n V_low
+ 817.000000n V_low
+ 817.000001n V_hig
+ 817.100000n V_hig
+ 817.100001n V_hig
+ 817.200000n V_hig
+ 817.200001n V_hig
+ 817.300000n V_hig
+ 817.300001n V_hig
+ 817.400000n V_hig
+ 817.400001n V_hig
+ 817.500000n V_hig
+ 817.500001n V_hig
+ 817.600000n V_hig
+ 817.600001n V_hig
+ 817.700000n V_hig
+ 817.700001n V_hig
+ 817.800000n V_hig
+ 817.800001n V_hig
+ 817.900000n V_hig
+ 817.900001n V_hig
+ 818.000000n V_hig
+ 818.000001n V_hig
+ 818.100000n V_hig
+ 818.100001n V_hig
+ 818.200000n V_hig
+ 818.200001n V_hig
+ 818.300000n V_hig
+ 818.300001n V_hig
+ 818.400000n V_hig
+ 818.400001n V_hig
+ 818.500000n V_hig
+ 818.500001n V_hig
+ 818.600000n V_hig
+ 818.600001n V_hig
+ 818.700000n V_hig
+ 818.700001n V_hig
+ 818.800000n V_hig
+ 818.800001n V_hig
+ 818.900000n V_hig
+ 818.900001n V_hig
+ 819.000000n V_hig
+ 819.000001n V_low
+ 819.100000n V_low
+ 819.100001n V_low
+ 819.200000n V_low
+ 819.200001n V_low
+ 819.300000n V_low
+ 819.300001n V_low
+ 819.400000n V_low
+ 819.400001n V_low
+ 819.500000n V_low
+ 819.500001n V_low
+ 819.600000n V_low
+ 819.600001n V_low
+ 819.700000n V_low
+ 819.700001n V_low
+ 819.800000n V_low
+ 819.800001n V_low
+ 819.900000n V_low
+ 819.900001n V_low
+ 820.000000n V_low
+ 820.000001n V_low
+ 820.100000n V_low
+ 820.100001n V_low
+ 820.200000n V_low
+ 820.200001n V_low
+ 820.300000n V_low
+ 820.300001n V_low
+ 820.400000n V_low
+ 820.400001n V_low
+ 820.500000n V_low
+ 820.500001n V_low
+ 820.600000n V_low
+ 820.600001n V_low
+ 820.700000n V_low
+ 820.700001n V_low
+ 820.800000n V_low
+ 820.800001n V_low
+ 820.900000n V_low
+ 820.900001n V_low
+ 821.000000n V_low
+ 821.000001n V_hig
+ 821.100000n V_hig
+ 821.100001n V_hig
+ 821.200000n V_hig
+ 821.200001n V_hig
+ 821.300000n V_hig
+ 821.300001n V_hig
+ 821.400000n V_hig
+ 821.400001n V_hig
+ 821.500000n V_hig
+ 821.500001n V_hig
+ 821.600000n V_hig
+ 821.600001n V_hig
+ 821.700000n V_hig
+ 821.700001n V_hig
+ 821.800000n V_hig
+ 821.800001n V_hig
+ 821.900000n V_hig
+ 821.900001n V_hig
+ 822.000000n V_hig
+ 822.000001n V_hig
+ 822.100000n V_hig
+ 822.100001n V_hig
+ 822.200000n V_hig
+ 822.200001n V_hig
+ 822.300000n V_hig
+ 822.300001n V_hig
+ 822.400000n V_hig
+ 822.400001n V_hig
+ 822.500000n V_hig
+ 822.500001n V_hig
+ 822.600000n V_hig
+ 822.600001n V_hig
+ 822.700000n V_hig
+ 822.700001n V_hig
+ 822.800000n V_hig
+ 822.800001n V_hig
+ 822.900000n V_hig
+ 822.900001n V_hig
+ 823.000000n V_hig
+ 823.000001n V_low
+ 823.100000n V_low
+ 823.100001n V_low
+ 823.200000n V_low
+ 823.200001n V_low
+ 823.300000n V_low
+ 823.300001n V_low
+ 823.400000n V_low
+ 823.400001n V_low
+ 823.500000n V_low
+ 823.500001n V_low
+ 823.600000n V_low
+ 823.600001n V_low
+ 823.700000n V_low
+ 823.700001n V_low
+ 823.800000n V_low
+ 823.800001n V_low
+ 823.900000n V_low
+ 823.900001n V_low
+ 824.000000n V_low
+ 824.000001n V_low
+ 824.100000n V_low
+ 824.100001n V_low
+ 824.200000n V_low
+ 824.200001n V_low
+ 824.300000n V_low
+ 824.300001n V_low
+ 824.400000n V_low
+ 824.400001n V_low
+ 824.500000n V_low
+ 824.500001n V_low
+ 824.600000n V_low
+ 824.600001n V_low
+ 824.700000n V_low
+ 824.700001n V_low
+ 824.800000n V_low
+ 824.800001n V_low
+ 824.900000n V_low
+ 824.900001n V_low
+ 825.000000n V_low
+ 825.000001n V_low
+ 825.100000n V_low
+ 825.100001n V_low
+ 825.200000n V_low
+ 825.200001n V_low
+ 825.300000n V_low
+ 825.300001n V_low
+ 825.400000n V_low
+ 825.400001n V_low
+ 825.500000n V_low
+ 825.500001n V_low
+ 825.600000n V_low
+ 825.600001n V_low
+ 825.700000n V_low
+ 825.700001n V_low
+ 825.800000n V_low
+ 825.800001n V_low
+ 825.900000n V_low
+ 825.900001n V_low
+ 826.000000n V_low
+ 826.000001n V_hig
+ 826.100000n V_hig
+ 826.100001n V_hig
+ 826.200000n V_hig
+ 826.200001n V_hig
+ 826.300000n V_hig
+ 826.300001n V_hig
+ 826.400000n V_hig
+ 826.400001n V_hig
+ 826.500000n V_hig
+ 826.500001n V_hig
+ 826.600000n V_hig
+ 826.600001n V_hig
+ 826.700000n V_hig
+ 826.700001n V_hig
+ 826.800000n V_hig
+ 826.800001n V_hig
+ 826.900000n V_hig
+ 826.900001n V_hig
+ 827.000000n V_hig
+ 827.000001n V_hig
+ 827.100000n V_hig
+ 827.100001n V_hig
+ 827.200000n V_hig
+ 827.200001n V_hig
+ 827.300000n V_hig
+ 827.300001n V_hig
+ 827.400000n V_hig
+ 827.400001n V_hig
+ 827.500000n V_hig
+ 827.500001n V_hig
+ 827.600000n V_hig
+ 827.600001n V_hig
+ 827.700000n V_hig
+ 827.700001n V_hig
+ 827.800000n V_hig
+ 827.800001n V_hig
+ 827.900000n V_hig
+ 827.900001n V_hig
+ 828.000000n V_hig
+ 828.000001n V_low
+ 828.100000n V_low
+ 828.100001n V_low
+ 828.200000n V_low
+ 828.200001n V_low
+ 828.300000n V_low
+ 828.300001n V_low
+ 828.400000n V_low
+ 828.400001n V_low
+ 828.500000n V_low
+ 828.500001n V_low
+ 828.600000n V_low
+ 828.600001n V_low
+ 828.700000n V_low
+ 828.700001n V_low
+ 828.800000n V_low
+ 828.800001n V_low
+ 828.900000n V_low
+ 828.900001n V_low
+ 829.000000n V_low
+ 829.000001n V_hig
+ 829.100000n V_hig
+ 829.100001n V_hig
+ 829.200000n V_hig
+ 829.200001n V_hig
+ 829.300000n V_hig
+ 829.300001n V_hig
+ 829.400000n V_hig
+ 829.400001n V_hig
+ 829.500000n V_hig
+ 829.500001n V_hig
+ 829.600000n V_hig
+ 829.600001n V_hig
+ 829.700000n V_hig
+ 829.700001n V_hig
+ 829.800000n V_hig
+ 829.800001n V_hig
+ 829.900000n V_hig
+ 829.900001n V_hig
+ 830.000000n V_hig
+ 830.000001n V_hig
+ 830.100000n V_hig
+ 830.100001n V_hig
+ 830.200000n V_hig
+ 830.200001n V_hig
+ 830.300000n V_hig
+ 830.300001n V_hig
+ 830.400000n V_hig
+ 830.400001n V_hig
+ 830.500000n V_hig
+ 830.500001n V_hig
+ 830.600000n V_hig
+ 830.600001n V_hig
+ 830.700000n V_hig
+ 830.700001n V_hig
+ 830.800000n V_hig
+ 830.800001n V_hig
+ 830.900000n V_hig
+ 830.900001n V_hig
+ 831.000000n V_hig
+ 831.000001n V_low
+ 831.100000n V_low
+ 831.100001n V_low
+ 831.200000n V_low
+ 831.200001n V_low
+ 831.300000n V_low
+ 831.300001n V_low
+ 831.400000n V_low
+ 831.400001n V_low
+ 831.500000n V_low
+ 831.500001n V_low
+ 831.600000n V_low
+ 831.600001n V_low
+ 831.700000n V_low
+ 831.700001n V_low
+ 831.800000n V_low
+ 831.800001n V_low
+ 831.900000n V_low
+ 831.900001n V_low
+ 832.000000n V_low
+ 832.000001n V_hig
+ 832.100000n V_hig
+ 832.100001n V_hig
+ 832.200000n V_hig
+ 832.200001n V_hig
+ 832.300000n V_hig
+ 832.300001n V_hig
+ 832.400000n V_hig
+ 832.400001n V_hig
+ 832.500000n V_hig
+ 832.500001n V_hig
+ 832.600000n V_hig
+ 832.600001n V_hig
+ 832.700000n V_hig
+ 832.700001n V_hig
+ 832.800000n V_hig
+ 832.800001n V_hig
+ 832.900000n V_hig
+ 832.900001n V_hig
+ 833.000000n V_hig
+ 833.000001n V_low
+ 833.100000n V_low
+ 833.100001n V_low
+ 833.200000n V_low
+ 833.200001n V_low
+ 833.300000n V_low
+ 833.300001n V_low
+ 833.400000n V_low
+ 833.400001n V_low
+ 833.500000n V_low
+ 833.500001n V_low
+ 833.600000n V_low
+ 833.600001n V_low
+ 833.700000n V_low
+ 833.700001n V_low
+ 833.800000n V_low
+ 833.800001n V_low
+ 833.900000n V_low
+ 833.900001n V_low
+ 834.000000n V_low
+ 834.000001n V_hig
+ 834.100000n V_hig
+ 834.100001n V_hig
+ 834.200000n V_hig
+ 834.200001n V_hig
+ 834.300000n V_hig
+ 834.300001n V_hig
+ 834.400000n V_hig
+ 834.400001n V_hig
+ 834.500000n V_hig
+ 834.500001n V_hig
+ 834.600000n V_hig
+ 834.600001n V_hig
+ 834.700000n V_hig
+ 834.700001n V_hig
+ 834.800000n V_hig
+ 834.800001n V_hig
+ 834.900000n V_hig
+ 834.900001n V_hig
+ 835.000000n V_hig
+ 835.000001n V_hig
+ 835.100000n V_hig
+ 835.100001n V_hig
+ 835.200000n V_hig
+ 835.200001n V_hig
+ 835.300000n V_hig
+ 835.300001n V_hig
+ 835.400000n V_hig
+ 835.400001n V_hig
+ 835.500000n V_hig
+ 835.500001n V_hig
+ 835.600000n V_hig
+ 835.600001n V_hig
+ 835.700000n V_hig
+ 835.700001n V_hig
+ 835.800000n V_hig
+ 835.800001n V_hig
+ 835.900000n V_hig
+ 835.900001n V_hig
+ 836.000000n V_hig
+ 836.000001n V_hig
+ 836.100000n V_hig
+ 836.100001n V_hig
+ 836.200000n V_hig
+ 836.200001n V_hig
+ 836.300000n V_hig
+ 836.300001n V_hig
+ 836.400000n V_hig
+ 836.400001n V_hig
+ 836.500000n V_hig
+ 836.500001n V_hig
+ 836.600000n V_hig
+ 836.600001n V_hig
+ 836.700000n V_hig
+ 836.700001n V_hig
+ 836.800000n V_hig
+ 836.800001n V_hig
+ 836.900000n V_hig
+ 836.900001n V_hig
+ 837.000000n V_hig
+ 837.000001n V_low
+ 837.100000n V_low
+ 837.100001n V_low
+ 837.200000n V_low
+ 837.200001n V_low
+ 837.300000n V_low
+ 837.300001n V_low
+ 837.400000n V_low
+ 837.400001n V_low
+ 837.500000n V_low
+ 837.500001n V_low
+ 837.600000n V_low
+ 837.600001n V_low
+ 837.700000n V_low
+ 837.700001n V_low
+ 837.800000n V_low
+ 837.800001n V_low
+ 837.900000n V_low
+ 837.900001n V_low
+ 838.000000n V_low
+ 838.000001n V_hig
+ 838.100000n V_hig
+ 838.100001n V_hig
+ 838.200000n V_hig
+ 838.200001n V_hig
+ 838.300000n V_hig
+ 838.300001n V_hig
+ 838.400000n V_hig
+ 838.400001n V_hig
+ 838.500000n V_hig
+ 838.500001n V_hig
+ 838.600000n V_hig
+ 838.600001n V_hig
+ 838.700000n V_hig
+ 838.700001n V_hig
+ 838.800000n V_hig
+ 838.800001n V_hig
+ 838.900000n V_hig
+ 838.900001n V_hig
+ 839.000000n V_hig
+ 839.000001n V_hig
+ 839.100000n V_hig
+ 839.100001n V_hig
+ 839.200000n V_hig
+ 839.200001n V_hig
+ 839.300000n V_hig
+ 839.300001n V_hig
+ 839.400000n V_hig
+ 839.400001n V_hig
+ 839.500000n V_hig
+ 839.500001n V_hig
+ 839.600000n V_hig
+ 839.600001n V_hig
+ 839.700000n V_hig
+ 839.700001n V_hig
+ 839.800000n V_hig
+ 839.800001n V_hig
+ 839.900000n V_hig
+ 839.900001n V_hig
+ 840.000000n V_hig
+ 840.000001n V_hig
+ 840.100000n V_hig
+ 840.100001n V_hig
+ 840.200000n V_hig
+ 840.200001n V_hig
+ 840.300000n V_hig
+ 840.300001n V_hig
+ 840.400000n V_hig
+ 840.400001n V_hig
+ 840.500000n V_hig
+ 840.500001n V_hig
+ 840.600000n V_hig
+ 840.600001n V_hig
+ 840.700000n V_hig
+ 840.700001n V_hig
+ 840.800000n V_hig
+ 840.800001n V_hig
+ 840.900000n V_hig
+ 840.900001n V_hig
+ 841.000000n V_hig
+ 841.000001n V_low
+ 841.100000n V_low
+ 841.100001n V_low
+ 841.200000n V_low
+ 841.200001n V_low
+ 841.300000n V_low
+ 841.300001n V_low
+ 841.400000n V_low
+ 841.400001n V_low
+ 841.500000n V_low
+ 841.500001n V_low
+ 841.600000n V_low
+ 841.600001n V_low
+ 841.700000n V_low
+ 841.700001n V_low
+ 841.800000n V_low
+ 841.800001n V_low
+ 841.900000n V_low
+ 841.900001n V_low
+ 842.000000n V_low
+ 842.000001n V_hig
+ 842.100000n V_hig
+ 842.100001n V_hig
+ 842.200000n V_hig
+ 842.200001n V_hig
+ 842.300000n V_hig
+ 842.300001n V_hig
+ 842.400000n V_hig
+ 842.400001n V_hig
+ 842.500000n V_hig
+ 842.500001n V_hig
+ 842.600000n V_hig
+ 842.600001n V_hig
+ 842.700000n V_hig
+ 842.700001n V_hig
+ 842.800000n V_hig
+ 842.800001n V_hig
+ 842.900000n V_hig
+ 842.900001n V_hig
+ 843.000000n V_hig
+ 843.000001n V_low
+ 843.100000n V_low
+ 843.100001n V_low
+ 843.200000n V_low
+ 843.200001n V_low
+ 843.300000n V_low
+ 843.300001n V_low
+ 843.400000n V_low
+ 843.400001n V_low
+ 843.500000n V_low
+ 843.500001n V_low
+ 843.600000n V_low
+ 843.600001n V_low
+ 843.700000n V_low
+ 843.700001n V_low
+ 843.800000n V_low
+ 843.800001n V_low
+ 843.900000n V_low
+ 843.900001n V_low
+ 844.000000n V_low
+ 844.000001n V_low
+ 844.100000n V_low
+ 844.100001n V_low
+ 844.200000n V_low
+ 844.200001n V_low
+ 844.300000n V_low
+ 844.300001n V_low
+ 844.400000n V_low
+ 844.400001n V_low
+ 844.500000n V_low
+ 844.500001n V_low
+ 844.600000n V_low
+ 844.600001n V_low
+ 844.700000n V_low
+ 844.700001n V_low
+ 844.800000n V_low
+ 844.800001n V_low
+ 844.900000n V_low
+ 844.900001n V_low
+ 845.000000n V_low
+ 845.000001n V_hig
+ 845.100000n V_hig
+ 845.100001n V_hig
+ 845.200000n V_hig
+ 845.200001n V_hig
+ 845.300000n V_hig
+ 845.300001n V_hig
+ 845.400000n V_hig
+ 845.400001n V_hig
+ 845.500000n V_hig
+ 845.500001n V_hig
+ 845.600000n V_hig
+ 845.600001n V_hig
+ 845.700000n V_hig
+ 845.700001n V_hig
+ 845.800000n V_hig
+ 845.800001n V_hig
+ 845.900000n V_hig
+ 845.900001n V_hig
+ 846.000000n V_hig
+ 846.000001n V_hig
+ 846.100000n V_hig
+ 846.100001n V_hig
+ 846.200000n V_hig
+ 846.200001n V_hig
+ 846.300000n V_hig
+ 846.300001n V_hig
+ 846.400000n V_hig
+ 846.400001n V_hig
+ 846.500000n V_hig
+ 846.500001n V_hig
+ 846.600000n V_hig
+ 846.600001n V_hig
+ 846.700000n V_hig
+ 846.700001n V_hig
+ 846.800000n V_hig
+ 846.800001n V_hig
+ 846.900000n V_hig
+ 846.900001n V_hig
+ 847.000000n V_hig
+ 847.000001n V_hig
+ 847.100000n V_hig
+ 847.100001n V_hig
+ 847.200000n V_hig
+ 847.200001n V_hig
+ 847.300000n V_hig
+ 847.300001n V_hig
+ 847.400000n V_hig
+ 847.400001n V_hig
+ 847.500000n V_hig
+ 847.500001n V_hig
+ 847.600000n V_hig
+ 847.600001n V_hig
+ 847.700000n V_hig
+ 847.700001n V_hig
+ 847.800000n V_hig
+ 847.800001n V_hig
+ 847.900000n V_hig
+ 847.900001n V_hig
+ 848.000000n V_hig
+ 848.000001n V_low
+ 848.100000n V_low
+ 848.100001n V_low
+ 848.200000n V_low
+ 848.200001n V_low
+ 848.300000n V_low
+ 848.300001n V_low
+ 848.400000n V_low
+ 848.400001n V_low
+ 848.500000n V_low
+ 848.500001n V_low
+ 848.600000n V_low
+ 848.600001n V_low
+ 848.700000n V_low
+ 848.700001n V_low
+ 848.800000n V_low
+ 848.800001n V_low
+ 848.900000n V_low
+ 848.900001n V_low
+ 849.000000n V_low
+ 849.000001n V_hig
+ 849.100000n V_hig
+ 849.100001n V_hig
+ 849.200000n V_hig
+ 849.200001n V_hig
+ 849.300000n V_hig
+ 849.300001n V_hig
+ 849.400000n V_hig
+ 849.400001n V_hig
+ 849.500000n V_hig
+ 849.500001n V_hig
+ 849.600000n V_hig
+ 849.600001n V_hig
+ 849.700000n V_hig
+ 849.700001n V_hig
+ 849.800000n V_hig
+ 849.800001n V_hig
+ 849.900000n V_hig
+ 849.900001n V_hig
+ 850.000000n V_hig
+ 850.000001n V_low
+ 850.100000n V_low
+ 850.100001n V_low
+ 850.200000n V_low
+ 850.200001n V_low
+ 850.300000n V_low
+ 850.300001n V_low
+ 850.400000n V_low
+ 850.400001n V_low
+ 850.500000n V_low
+ 850.500001n V_low
+ 850.600000n V_low
+ 850.600001n V_low
+ 850.700000n V_low
+ 850.700001n V_low
+ 850.800000n V_low
+ 850.800001n V_low
+ 850.900000n V_low
+ 850.900001n V_low
+ 851.000000n V_low
+ 851.000001n V_hig
+ 851.100000n V_hig
+ 851.100001n V_hig
+ 851.200000n V_hig
+ 851.200001n V_hig
+ 851.300000n V_hig
+ 851.300001n V_hig
+ 851.400000n V_hig
+ 851.400001n V_hig
+ 851.500000n V_hig
+ 851.500001n V_hig
+ 851.600000n V_hig
+ 851.600001n V_hig
+ 851.700000n V_hig
+ 851.700001n V_hig
+ 851.800000n V_hig
+ 851.800001n V_hig
+ 851.900000n V_hig
+ 851.900001n V_hig
+ 852.000000n V_hig
+ 852.000001n V_hig
+ 852.100000n V_hig
+ 852.100001n V_hig
+ 852.200000n V_hig
+ 852.200001n V_hig
+ 852.300000n V_hig
+ 852.300001n V_hig
+ 852.400000n V_hig
+ 852.400001n V_hig
+ 852.500000n V_hig
+ 852.500001n V_hig
+ 852.600000n V_hig
+ 852.600001n V_hig
+ 852.700000n V_hig
+ 852.700001n V_hig
+ 852.800000n V_hig
+ 852.800001n V_hig
+ 852.900000n V_hig
+ 852.900001n V_hig
+ 853.000000n V_hig
+ 853.000001n V_low
+ 853.100000n V_low
+ 853.100001n V_low
+ 853.200000n V_low
+ 853.200001n V_low
+ 853.300000n V_low
+ 853.300001n V_low
+ 853.400000n V_low
+ 853.400001n V_low
+ 853.500000n V_low
+ 853.500001n V_low
+ 853.600000n V_low
+ 853.600001n V_low
+ 853.700000n V_low
+ 853.700001n V_low
+ 853.800000n V_low
+ 853.800001n V_low
+ 853.900000n V_low
+ 853.900001n V_low
+ 854.000000n V_low
+ 854.000001n V_hig
+ 854.100000n V_hig
+ 854.100001n V_hig
+ 854.200000n V_hig
+ 854.200001n V_hig
+ 854.300000n V_hig
+ 854.300001n V_hig
+ 854.400000n V_hig
+ 854.400001n V_hig
+ 854.500000n V_hig
+ 854.500001n V_hig
+ 854.600000n V_hig
+ 854.600001n V_hig
+ 854.700000n V_hig
+ 854.700001n V_hig
+ 854.800000n V_hig
+ 854.800001n V_hig
+ 854.900000n V_hig
+ 854.900001n V_hig
+ 855.000000n V_hig
+ 855.000001n V_low
+ 855.100000n V_low
+ 855.100001n V_low
+ 855.200000n V_low
+ 855.200001n V_low
+ 855.300000n V_low
+ 855.300001n V_low
+ 855.400000n V_low
+ 855.400001n V_low
+ 855.500000n V_low
+ 855.500001n V_low
+ 855.600000n V_low
+ 855.600001n V_low
+ 855.700000n V_low
+ 855.700001n V_low
+ 855.800000n V_low
+ 855.800001n V_low
+ 855.900000n V_low
+ 855.900001n V_low
+ 856.000000n V_low
+ 856.000001n V_low
+ 856.100000n V_low
+ 856.100001n V_low
+ 856.200000n V_low
+ 856.200001n V_low
+ 856.300000n V_low
+ 856.300001n V_low
+ 856.400000n V_low
+ 856.400001n V_low
+ 856.500000n V_low
+ 856.500001n V_low
+ 856.600000n V_low
+ 856.600001n V_low
+ 856.700000n V_low
+ 856.700001n V_low
+ 856.800000n V_low
+ 856.800001n V_low
+ 856.900000n V_low
+ 856.900001n V_low
+ 857.000000n V_low
+ 857.000001n V_hig
+ 857.100000n V_hig
+ 857.100001n V_hig
+ 857.200000n V_hig
+ 857.200001n V_hig
+ 857.300000n V_hig
+ 857.300001n V_hig
+ 857.400000n V_hig
+ 857.400001n V_hig
+ 857.500000n V_hig
+ 857.500001n V_hig
+ 857.600000n V_hig
+ 857.600001n V_hig
+ 857.700000n V_hig
+ 857.700001n V_hig
+ 857.800000n V_hig
+ 857.800001n V_hig
+ 857.900000n V_hig
+ 857.900001n V_hig
+ 858.000000n V_hig
+ 858.000001n V_low
+ 858.100000n V_low
+ 858.100001n V_low
+ 858.200000n V_low
+ 858.200001n V_low
+ 858.300000n V_low
+ 858.300001n V_low
+ 858.400000n V_low
+ 858.400001n V_low
+ 858.500000n V_low
+ 858.500001n V_low
+ 858.600000n V_low
+ 858.600001n V_low
+ 858.700000n V_low
+ 858.700001n V_low
+ 858.800000n V_low
+ 858.800001n V_low
+ 858.900000n V_low
+ 858.900001n V_low
+ 859.000000n V_low
+ 859.000001n V_hig
+ 859.100000n V_hig
+ 859.100001n V_hig
+ 859.200000n V_hig
+ 859.200001n V_hig
+ 859.300000n V_hig
+ 859.300001n V_hig
+ 859.400000n V_hig
+ 859.400001n V_hig
+ 859.500000n V_hig
+ 859.500001n V_hig
+ 859.600000n V_hig
+ 859.600001n V_hig
+ 859.700000n V_hig
+ 859.700001n V_hig
+ 859.800000n V_hig
+ 859.800001n V_hig
+ 859.900000n V_hig
+ 859.900001n V_hig
+ 860.000000n V_hig
+ 860.000001n V_low
+ 860.100000n V_low
+ 860.100001n V_low
+ 860.200000n V_low
+ 860.200001n V_low
+ 860.300000n V_low
+ 860.300001n V_low
+ 860.400000n V_low
+ 860.400001n V_low
+ 860.500000n V_low
+ 860.500001n V_low
+ 860.600000n V_low
+ 860.600001n V_low
+ 860.700000n V_low
+ 860.700001n V_low
+ 860.800000n V_low
+ 860.800001n V_low
+ 860.900000n V_low
+ 860.900001n V_low
+ 861.000000n V_low
+ 861.000001n V_low
+ 861.100000n V_low
+ 861.100001n V_low
+ 861.200000n V_low
+ 861.200001n V_low
+ 861.300000n V_low
+ 861.300001n V_low
+ 861.400000n V_low
+ 861.400001n V_low
+ 861.500000n V_low
+ 861.500001n V_low
+ 861.600000n V_low
+ 861.600001n V_low
+ 861.700000n V_low
+ 861.700001n V_low
+ 861.800000n V_low
+ 861.800001n V_low
+ 861.900000n V_low
+ 861.900001n V_low
+ 862.000000n V_low
+ 862.000001n V_hig
+ 862.100000n V_hig
+ 862.100001n V_hig
+ 862.200000n V_hig
+ 862.200001n V_hig
+ 862.300000n V_hig
+ 862.300001n V_hig
+ 862.400000n V_hig
+ 862.400001n V_hig
+ 862.500000n V_hig
+ 862.500001n V_hig
+ 862.600000n V_hig
+ 862.600001n V_hig
+ 862.700000n V_hig
+ 862.700001n V_hig
+ 862.800000n V_hig
+ 862.800001n V_hig
+ 862.900000n V_hig
+ 862.900001n V_hig
+ 863.000000n V_hig
+ 863.000001n V_hig
+ 863.100000n V_hig
+ 863.100001n V_hig
+ 863.200000n V_hig
+ 863.200001n V_hig
+ 863.300000n V_hig
+ 863.300001n V_hig
+ 863.400000n V_hig
+ 863.400001n V_hig
+ 863.500000n V_hig
+ 863.500001n V_hig
+ 863.600000n V_hig
+ 863.600001n V_hig
+ 863.700000n V_hig
+ 863.700001n V_hig
+ 863.800000n V_hig
+ 863.800001n V_hig
+ 863.900000n V_hig
+ 863.900001n V_hig
+ 864.000000n V_hig
+ 864.000001n V_low
+ 864.100000n V_low
+ 864.100001n V_low
+ 864.200000n V_low
+ 864.200001n V_low
+ 864.300000n V_low
+ 864.300001n V_low
+ 864.400000n V_low
+ 864.400001n V_low
+ 864.500000n V_low
+ 864.500001n V_low
+ 864.600000n V_low
+ 864.600001n V_low
+ 864.700000n V_low
+ 864.700001n V_low
+ 864.800000n V_low
+ 864.800001n V_low
+ 864.900000n V_low
+ 864.900001n V_low
+ 865.000000n V_low
+ 865.000001n V_low
+ 865.100000n V_low
+ 865.100001n V_low
+ 865.200000n V_low
+ 865.200001n V_low
+ 865.300000n V_low
+ 865.300001n V_low
+ 865.400000n V_low
+ 865.400001n V_low
+ 865.500000n V_low
+ 865.500001n V_low
+ 865.600000n V_low
+ 865.600001n V_low
+ 865.700000n V_low
+ 865.700001n V_low
+ 865.800000n V_low
+ 865.800001n V_low
+ 865.900000n V_low
+ 865.900001n V_low
+ 866.000000n V_low
+ 866.000001n V_low
+ 866.100000n V_low
+ 866.100001n V_low
+ 866.200000n V_low
+ 866.200001n V_low
+ 866.300000n V_low
+ 866.300001n V_low
+ 866.400000n V_low
+ 866.400001n V_low
+ 866.500000n V_low
+ 866.500001n V_low
+ 866.600000n V_low
+ 866.600001n V_low
+ 866.700000n V_low
+ 866.700001n V_low
+ 866.800000n V_low
+ 866.800001n V_low
+ 866.900000n V_low
+ 866.900001n V_low
+ 867.000000n V_low
+ 867.000001n V_low
+ 867.100000n V_low
+ 867.100001n V_low
+ 867.200000n V_low
+ 867.200001n V_low
+ 867.300000n V_low
+ 867.300001n V_low
+ 867.400000n V_low
+ 867.400001n V_low
+ 867.500000n V_low
+ 867.500001n V_low
+ 867.600000n V_low
+ 867.600001n V_low
+ 867.700000n V_low
+ 867.700001n V_low
+ 867.800000n V_low
+ 867.800001n V_low
+ 867.900000n V_low
+ 867.900001n V_low
+ 868.000000n V_low
+ 868.000001n V_hig
+ 868.100000n V_hig
+ 868.100001n V_hig
+ 868.200000n V_hig
+ 868.200001n V_hig
+ 868.300000n V_hig
+ 868.300001n V_hig
+ 868.400000n V_hig
+ 868.400001n V_hig
+ 868.500000n V_hig
+ 868.500001n V_hig
+ 868.600000n V_hig
+ 868.600001n V_hig
+ 868.700000n V_hig
+ 868.700001n V_hig
+ 868.800000n V_hig
+ 868.800001n V_hig
+ 868.900000n V_hig
+ 868.900001n V_hig
+ 869.000000n V_hig
+ 869.000001n V_hig
+ 869.100000n V_hig
+ 869.100001n V_hig
+ 869.200000n V_hig
+ 869.200001n V_hig
+ 869.300000n V_hig
+ 869.300001n V_hig
+ 869.400000n V_hig
+ 869.400001n V_hig
+ 869.500000n V_hig
+ 869.500001n V_hig
+ 869.600000n V_hig
+ 869.600001n V_hig
+ 869.700000n V_hig
+ 869.700001n V_hig
+ 869.800000n V_hig
+ 869.800001n V_hig
+ 869.900000n V_hig
+ 869.900001n V_hig
+ 870.000000n V_hig
+ 870.000001n V_low
+ 870.100000n V_low
+ 870.100001n V_low
+ 870.200000n V_low
+ 870.200001n V_low
+ 870.300000n V_low
+ 870.300001n V_low
+ 870.400000n V_low
+ 870.400001n V_low
+ 870.500000n V_low
+ 870.500001n V_low
+ 870.600000n V_low
+ 870.600001n V_low
+ 870.700000n V_low
+ 870.700001n V_low
+ 870.800000n V_low
+ 870.800001n V_low
+ 870.900000n V_low
+ 870.900001n V_low
+ 871.000000n V_low
+ 871.000001n V_low
+ 871.100000n V_low
+ 871.100001n V_low
+ 871.200000n V_low
+ 871.200001n V_low
+ 871.300000n V_low
+ 871.300001n V_low
+ 871.400000n V_low
+ 871.400001n V_low
+ 871.500000n V_low
+ 871.500001n V_low
+ 871.600000n V_low
+ 871.600001n V_low
+ 871.700000n V_low
+ 871.700001n V_low
+ 871.800000n V_low
+ 871.800001n V_low
+ 871.900000n V_low
+ 871.900001n V_low
+ 872.000000n V_low
+ 872.000001n V_hig
+ 872.100000n V_hig
+ 872.100001n V_hig
+ 872.200000n V_hig
+ 872.200001n V_hig
+ 872.300000n V_hig
+ 872.300001n V_hig
+ 872.400000n V_hig
+ 872.400001n V_hig
+ 872.500000n V_hig
+ 872.500001n V_hig
+ 872.600000n V_hig
+ 872.600001n V_hig
+ 872.700000n V_hig
+ 872.700001n V_hig
+ 872.800000n V_hig
+ 872.800001n V_hig
+ 872.900000n V_hig
+ 872.900001n V_hig
+ 873.000000n V_hig
+ 873.000001n V_hig
+ 873.100000n V_hig
+ 873.100001n V_hig
+ 873.200000n V_hig
+ 873.200001n V_hig
+ 873.300000n V_hig
+ 873.300001n V_hig
+ 873.400000n V_hig
+ 873.400001n V_hig
+ 873.500000n V_hig
+ 873.500001n V_hig
+ 873.600000n V_hig
+ 873.600001n V_hig
+ 873.700000n V_hig
+ 873.700001n V_hig
+ 873.800000n V_hig
+ 873.800001n V_hig
+ 873.900000n V_hig
+ 873.900001n V_hig
+ 874.000000n V_hig
+ 874.000001n V_low
+ 874.100000n V_low
+ 874.100001n V_low
+ 874.200000n V_low
+ 874.200001n V_low
+ 874.300000n V_low
+ 874.300001n V_low
+ 874.400000n V_low
+ 874.400001n V_low
+ 874.500000n V_low
+ 874.500001n V_low
+ 874.600000n V_low
+ 874.600001n V_low
+ 874.700000n V_low
+ 874.700001n V_low
+ 874.800000n V_low
+ 874.800001n V_low
+ 874.900000n V_low
+ 874.900001n V_low
+ 875.000000n V_low
+ 875.000001n V_low
+ 875.100000n V_low
+ 875.100001n V_low
+ 875.200000n V_low
+ 875.200001n V_low
+ 875.300000n V_low
+ 875.300001n V_low
+ 875.400000n V_low
+ 875.400001n V_low
+ 875.500000n V_low
+ 875.500001n V_low
+ 875.600000n V_low
+ 875.600001n V_low
+ 875.700000n V_low
+ 875.700001n V_low
+ 875.800000n V_low
+ 875.800001n V_low
+ 875.900000n V_low
+ 875.900001n V_low
+ 876.000000n V_low
+ 876.000001n V_hig
+ 876.100000n V_hig
+ 876.100001n V_hig
+ 876.200000n V_hig
+ 876.200001n V_hig
+ 876.300000n V_hig
+ 876.300001n V_hig
+ 876.400000n V_hig
+ 876.400001n V_hig
+ 876.500000n V_hig
+ 876.500001n V_hig
+ 876.600000n V_hig
+ 876.600001n V_hig
+ 876.700000n V_hig
+ 876.700001n V_hig
+ 876.800000n V_hig
+ 876.800001n V_hig
+ 876.900000n V_hig
+ 876.900001n V_hig
+ 877.000000n V_hig
+ 877.000001n V_hig
+ 877.100000n V_hig
+ 877.100001n V_hig
+ 877.200000n V_hig
+ 877.200001n V_hig
+ 877.300000n V_hig
+ 877.300001n V_hig
+ 877.400000n V_hig
+ 877.400001n V_hig
+ 877.500000n V_hig
+ 877.500001n V_hig
+ 877.600000n V_hig
+ 877.600001n V_hig
+ 877.700000n V_hig
+ 877.700001n V_hig
+ 877.800000n V_hig
+ 877.800001n V_hig
+ 877.900000n V_hig
+ 877.900001n V_hig
+ 878.000000n V_hig
+ 878.000001n V_low
+ 878.100000n V_low
+ 878.100001n V_low
+ 878.200000n V_low
+ 878.200001n V_low
+ 878.300000n V_low
+ 878.300001n V_low
+ 878.400000n V_low
+ 878.400001n V_low
+ 878.500000n V_low
+ 878.500001n V_low
+ 878.600000n V_low
+ 878.600001n V_low
+ 878.700000n V_low
+ 878.700001n V_low
+ 878.800000n V_low
+ 878.800001n V_low
+ 878.900000n V_low
+ 878.900001n V_low
+ 879.000000n V_low
+ 879.000001n V_low
+ 879.100000n V_low
+ 879.100001n V_low
+ 879.200000n V_low
+ 879.200001n V_low
+ 879.300000n V_low
+ 879.300001n V_low
+ 879.400000n V_low
+ 879.400001n V_low
+ 879.500000n V_low
+ 879.500001n V_low
+ 879.600000n V_low
+ 879.600001n V_low
+ 879.700000n V_low
+ 879.700001n V_low
+ 879.800000n V_low
+ 879.800001n V_low
+ 879.900000n V_low
+ 879.900001n V_low
+ 880.000000n V_low
+ 880.000001n V_low
+ 880.100000n V_low
+ 880.100001n V_low
+ 880.200000n V_low
+ 880.200001n V_low
+ 880.300000n V_low
+ 880.300001n V_low
+ 880.400000n V_low
+ 880.400001n V_low
+ 880.500000n V_low
+ 880.500001n V_low
+ 880.600000n V_low
+ 880.600001n V_low
+ 880.700000n V_low
+ 880.700001n V_low
+ 880.800000n V_low
+ 880.800001n V_low
+ 880.900000n V_low
+ 880.900001n V_low
+ 881.000000n V_low
+ 881.000001n V_low
+ 881.100000n V_low
+ 881.100001n V_low
+ 881.200000n V_low
+ 881.200001n V_low
+ 881.300000n V_low
+ 881.300001n V_low
+ 881.400000n V_low
+ 881.400001n V_low
+ 881.500000n V_low
+ 881.500001n V_low
+ 881.600000n V_low
+ 881.600001n V_low
+ 881.700000n V_low
+ 881.700001n V_low
+ 881.800000n V_low
+ 881.800001n V_low
+ 881.900000n V_low
+ 881.900001n V_low
+ 882.000000n V_low
+ 882.000001n V_low
+ 882.100000n V_low
+ 882.100001n V_low
+ 882.200000n V_low
+ 882.200001n V_low
+ 882.300000n V_low
+ 882.300001n V_low
+ 882.400000n V_low
+ 882.400001n V_low
+ 882.500000n V_low
+ 882.500001n V_low
+ 882.600000n V_low
+ 882.600001n V_low
+ 882.700000n V_low
+ 882.700001n V_low
+ 882.800000n V_low
+ 882.800001n V_low
+ 882.900000n V_low
+ 882.900001n V_low
+ 883.000000n V_low
+ 883.000001n V_hig
+ 883.100000n V_hig
+ 883.100001n V_hig
+ 883.200000n V_hig
+ 883.200001n V_hig
+ 883.300000n V_hig
+ 883.300001n V_hig
+ 883.400000n V_hig
+ 883.400001n V_hig
+ 883.500000n V_hig
+ 883.500001n V_hig
+ 883.600000n V_hig
+ 883.600001n V_hig
+ 883.700000n V_hig
+ 883.700001n V_hig
+ 883.800000n V_hig
+ 883.800001n V_hig
+ 883.900000n V_hig
+ 883.900001n V_hig
+ 884.000000n V_hig
+ 884.000001n V_hig
+ 884.100000n V_hig
+ 884.100001n V_hig
+ 884.200000n V_hig
+ 884.200001n V_hig
+ 884.300000n V_hig
+ 884.300001n V_hig
+ 884.400000n V_hig
+ 884.400001n V_hig
+ 884.500000n V_hig
+ 884.500001n V_hig
+ 884.600000n V_hig
+ 884.600001n V_hig
+ 884.700000n V_hig
+ 884.700001n V_hig
+ 884.800000n V_hig
+ 884.800001n V_hig
+ 884.900000n V_hig
+ 884.900001n V_hig
+ 885.000000n V_hig
+ 885.000001n V_hig
+ 885.100000n V_hig
+ 885.100001n V_hig
+ 885.200000n V_hig
+ 885.200001n V_hig
+ 885.300000n V_hig
+ 885.300001n V_hig
+ 885.400000n V_hig
+ 885.400001n V_hig
+ 885.500000n V_hig
+ 885.500001n V_hig
+ 885.600000n V_hig
+ 885.600001n V_hig
+ 885.700000n V_hig
+ 885.700001n V_hig
+ 885.800000n V_hig
+ 885.800001n V_hig
+ 885.900000n V_hig
+ 885.900001n V_hig
+ 886.000000n V_hig
+ 886.000001n V_low
+ 886.100000n V_low
+ 886.100001n V_low
+ 886.200000n V_low
+ 886.200001n V_low
+ 886.300000n V_low
+ 886.300001n V_low
+ 886.400000n V_low
+ 886.400001n V_low
+ 886.500000n V_low
+ 886.500001n V_low
+ 886.600000n V_low
+ 886.600001n V_low
+ 886.700000n V_low
+ 886.700001n V_low
+ 886.800000n V_low
+ 886.800001n V_low
+ 886.900000n V_low
+ 886.900001n V_low
+ 887.000000n V_low
+ 887.000001n V_hig
+ 887.100000n V_hig
+ 887.100001n V_hig
+ 887.200000n V_hig
+ 887.200001n V_hig
+ 887.300000n V_hig
+ 887.300001n V_hig
+ 887.400000n V_hig
+ 887.400001n V_hig
+ 887.500000n V_hig
+ 887.500001n V_hig
+ 887.600000n V_hig
+ 887.600001n V_hig
+ 887.700000n V_hig
+ 887.700001n V_hig
+ 887.800000n V_hig
+ 887.800001n V_hig
+ 887.900000n V_hig
+ 887.900001n V_hig
+ 888.000000n V_hig
+ 888.000001n V_hig
+ 888.100000n V_hig
+ 888.100001n V_hig
+ 888.200000n V_hig
+ 888.200001n V_hig
+ 888.300000n V_hig
+ 888.300001n V_hig
+ 888.400000n V_hig
+ 888.400001n V_hig
+ 888.500000n V_hig
+ 888.500001n V_hig
+ 888.600000n V_hig
+ 888.600001n V_hig
+ 888.700000n V_hig
+ 888.700001n V_hig
+ 888.800000n V_hig
+ 888.800001n V_hig
+ 888.900000n V_hig
+ 888.900001n V_hig
+ 889.000000n V_hig
+ 889.000001n V_low
+ 889.100000n V_low
+ 889.100001n V_low
+ 889.200000n V_low
+ 889.200001n V_low
+ 889.300000n V_low
+ 889.300001n V_low
+ 889.400000n V_low
+ 889.400001n V_low
+ 889.500000n V_low
+ 889.500001n V_low
+ 889.600000n V_low
+ 889.600001n V_low
+ 889.700000n V_low
+ 889.700001n V_low
+ 889.800000n V_low
+ 889.800001n V_low
+ 889.900000n V_low
+ 889.900001n V_low
+ 890.000000n V_low
+ 890.000001n V_low
+ 890.100000n V_low
+ 890.100001n V_low
+ 890.200000n V_low
+ 890.200001n V_low
+ 890.300000n V_low
+ 890.300001n V_low
+ 890.400000n V_low
+ 890.400001n V_low
+ 890.500000n V_low
+ 890.500001n V_low
+ 890.600000n V_low
+ 890.600001n V_low
+ 890.700000n V_low
+ 890.700001n V_low
+ 890.800000n V_low
+ 890.800001n V_low
+ 890.900000n V_low
+ 890.900001n V_low
+ 891.000000n V_low
+ 891.000001n V_hig
+ 891.100000n V_hig
+ 891.100001n V_hig
+ 891.200000n V_hig
+ 891.200001n V_hig
+ 891.300000n V_hig
+ 891.300001n V_hig
+ 891.400000n V_hig
+ 891.400001n V_hig
+ 891.500000n V_hig
+ 891.500001n V_hig
+ 891.600000n V_hig
+ 891.600001n V_hig
+ 891.700000n V_hig
+ 891.700001n V_hig
+ 891.800000n V_hig
+ 891.800001n V_hig
+ 891.900000n V_hig
+ 891.900001n V_hig
+ 892.000000n V_hig
+ 892.000001n V_hig
+ 892.100000n V_hig
+ 892.100001n V_hig
+ 892.200000n V_hig
+ 892.200001n V_hig
+ 892.300000n V_hig
+ 892.300001n V_hig
+ 892.400000n V_hig
+ 892.400001n V_hig
+ 892.500000n V_hig
+ 892.500001n V_hig
+ 892.600000n V_hig
+ 892.600001n V_hig
+ 892.700000n V_hig
+ 892.700001n V_hig
+ 892.800000n V_hig
+ 892.800001n V_hig
+ 892.900000n V_hig
+ 892.900001n V_hig
+ 893.000000n V_hig
+ 893.000001n V_hig
+ 893.100000n V_hig
+ 893.100001n V_hig
+ 893.200000n V_hig
+ 893.200001n V_hig
+ 893.300000n V_hig
+ 893.300001n V_hig
+ 893.400000n V_hig
+ 893.400001n V_hig
+ 893.500000n V_hig
+ 893.500001n V_hig
+ 893.600000n V_hig
+ 893.600001n V_hig
+ 893.700000n V_hig
+ 893.700001n V_hig
+ 893.800000n V_hig
+ 893.800001n V_hig
+ 893.900000n V_hig
+ 893.900001n V_hig
+ 894.000000n V_hig
+ 894.000001n V_low
+ 894.100000n V_low
+ 894.100001n V_low
+ 894.200000n V_low
+ 894.200001n V_low
+ 894.300000n V_low
+ 894.300001n V_low
+ 894.400000n V_low
+ 894.400001n V_low
+ 894.500000n V_low
+ 894.500001n V_low
+ 894.600000n V_low
+ 894.600001n V_low
+ 894.700000n V_low
+ 894.700001n V_low
+ 894.800000n V_low
+ 894.800001n V_low
+ 894.900000n V_low
+ 894.900001n V_low
+ 895.000000n V_low
+ 895.000001n V_hig
+ 895.100000n V_hig
+ 895.100001n V_hig
+ 895.200000n V_hig
+ 895.200001n V_hig
+ 895.300000n V_hig
+ 895.300001n V_hig
+ 895.400000n V_hig
+ 895.400001n V_hig
+ 895.500000n V_hig
+ 895.500001n V_hig
+ 895.600000n V_hig
+ 895.600001n V_hig
+ 895.700000n V_hig
+ 895.700001n V_hig
+ 895.800000n V_hig
+ 895.800001n V_hig
+ 895.900000n V_hig
+ 895.900001n V_hig
+ 896.000000n V_hig
+ 896.000001n V_hig
+ 896.100000n V_hig
+ 896.100001n V_hig
+ 896.200000n V_hig
+ 896.200001n V_hig
+ 896.300000n V_hig
+ 896.300001n V_hig
+ 896.400000n V_hig
+ 896.400001n V_hig
+ 896.500000n V_hig
+ 896.500001n V_hig
+ 896.600000n V_hig
+ 896.600001n V_hig
+ 896.700000n V_hig
+ 896.700001n V_hig
+ 896.800000n V_hig
+ 896.800001n V_hig
+ 896.900000n V_hig
+ 896.900001n V_hig
+ 897.000000n V_hig
+ 897.000001n V_hig
+ 897.100000n V_hig
+ 897.100001n V_hig
+ 897.200000n V_hig
+ 897.200001n V_hig
+ 897.300000n V_hig
+ 897.300001n V_hig
+ 897.400000n V_hig
+ 897.400001n V_hig
+ 897.500000n V_hig
+ 897.500001n V_hig
+ 897.600000n V_hig
+ 897.600001n V_hig
+ 897.700000n V_hig
+ 897.700001n V_hig
+ 897.800000n V_hig
+ 897.800001n V_hig
+ 897.900000n V_hig
+ 897.900001n V_hig
+ 898.000000n V_hig
+ 898.000001n V_low
+ 898.100000n V_low
+ 898.100001n V_low
+ 898.200000n V_low
+ 898.200001n V_low
+ 898.300000n V_low
+ 898.300001n V_low
+ 898.400000n V_low
+ 898.400001n V_low
+ 898.500000n V_low
+ 898.500001n V_low
+ 898.600000n V_low
+ 898.600001n V_low
+ 898.700000n V_low
+ 898.700001n V_low
+ 898.800000n V_low
+ 898.800001n V_low
+ 898.900000n V_low
+ 898.900001n V_low
+ 899.000000n V_low
+ 899.000001n V_low
+ 899.100000n V_low
+ 899.100001n V_low
+ 899.200000n V_low
+ 899.200001n V_low
+ 899.300000n V_low
+ 899.300001n V_low
+ 899.400000n V_low
+ 899.400001n V_low
+ 899.500000n V_low
+ 899.500001n V_low
+ 899.600000n V_low
+ 899.600001n V_low
+ 899.700000n V_low
+ 899.700001n V_low
+ 899.800000n V_low
+ 899.800001n V_low
+ 899.900000n V_low
+ 899.900001n V_low
+ 900.000000n V_low
+ 900.000001n V_hig
+ 900.100000n V_hig
+ 900.100001n V_hig
+ 900.200000n V_hig
+ 900.200001n V_hig
+ 900.300000n V_hig
+ 900.300001n V_hig
+ 900.400000n V_hig
+ 900.400001n V_hig
+ 900.500000n V_hig
+ 900.500001n V_hig
+ 900.600000n V_hig
+ 900.600001n V_hig
+ 900.700000n V_hig
+ 900.700001n V_hig
+ 900.800000n V_hig
+ 900.800001n V_hig
+ 900.900000n V_hig
+ 900.900001n V_hig
+ 901.000000n V_hig
+ 901.000001n V_hig
+ 901.100000n V_hig
+ 901.100001n V_hig
+ 901.200000n V_hig
+ 901.200001n V_hig
+ 901.300000n V_hig
+ 901.300001n V_hig
+ 901.400000n V_hig
+ 901.400001n V_hig
+ 901.500000n V_hig
+ 901.500001n V_hig
+ 901.600000n V_hig
+ 901.600001n V_hig
+ 901.700000n V_hig
+ 901.700001n V_hig
+ 901.800000n V_hig
+ 901.800001n V_hig
+ 901.900000n V_hig
+ 901.900001n V_hig
+ 902.000000n V_hig
+ 902.000001n V_hig
+ 902.100000n V_hig
+ 902.100001n V_hig
+ 902.200000n V_hig
+ 902.200001n V_hig
+ 902.300000n V_hig
+ 902.300001n V_hig
+ 902.400000n V_hig
+ 902.400001n V_hig
+ 902.500000n V_hig
+ 902.500001n V_hig
+ 902.600000n V_hig
+ 902.600001n V_hig
+ 902.700000n V_hig
+ 902.700001n V_hig
+ 902.800000n V_hig
+ 902.800001n V_hig
+ 902.900000n V_hig
+ 902.900001n V_hig
+ 903.000000n V_hig
+ 903.000001n V_low
+ 903.100000n V_low
+ 903.100001n V_low
+ 903.200000n V_low
+ 903.200001n V_low
+ 903.300000n V_low
+ 903.300001n V_low
+ 903.400000n V_low
+ 903.400001n V_low
+ 903.500000n V_low
+ 903.500001n V_low
+ 903.600000n V_low
+ 903.600001n V_low
+ 903.700000n V_low
+ 903.700001n V_low
+ 903.800000n V_low
+ 903.800001n V_low
+ 903.900000n V_low
+ 903.900001n V_low
+ 904.000000n V_low
+ 904.000001n V_hig
+ 904.100000n V_hig
+ 904.100001n V_hig
+ 904.200000n V_hig
+ 904.200001n V_hig
+ 904.300000n V_hig
+ 904.300001n V_hig
+ 904.400000n V_hig
+ 904.400001n V_hig
+ 904.500000n V_hig
+ 904.500001n V_hig
+ 904.600000n V_hig
+ 904.600001n V_hig
+ 904.700000n V_hig
+ 904.700001n V_hig
+ 904.800000n V_hig
+ 904.800001n V_hig
+ 904.900000n V_hig
+ 904.900001n V_hig
+ 905.000000n V_hig
+ 905.000001n V_hig
+ 905.100000n V_hig
+ 905.100001n V_hig
+ 905.200000n V_hig
+ 905.200001n V_hig
+ 905.300000n V_hig
+ 905.300001n V_hig
+ 905.400000n V_hig
+ 905.400001n V_hig
+ 905.500000n V_hig
+ 905.500001n V_hig
+ 905.600000n V_hig
+ 905.600001n V_hig
+ 905.700000n V_hig
+ 905.700001n V_hig
+ 905.800000n V_hig
+ 905.800001n V_hig
+ 905.900000n V_hig
+ 905.900001n V_hig
+ 906.000000n V_hig
+ 906.000001n V_low
+ 906.100000n V_low
+ 906.100001n V_low
+ 906.200000n V_low
+ 906.200001n V_low
+ 906.300000n V_low
+ 906.300001n V_low
+ 906.400000n V_low
+ 906.400001n V_low
+ 906.500000n V_low
+ 906.500001n V_low
+ 906.600000n V_low
+ 906.600001n V_low
+ 906.700000n V_low
+ 906.700001n V_low
+ 906.800000n V_low
+ 906.800001n V_low
+ 906.900000n V_low
+ 906.900001n V_low
+ 907.000000n V_low
+ 907.000001n V_low
+ 907.100000n V_low
+ 907.100001n V_low
+ 907.200000n V_low
+ 907.200001n V_low
+ 907.300000n V_low
+ 907.300001n V_low
+ 907.400000n V_low
+ 907.400001n V_low
+ 907.500000n V_low
+ 907.500001n V_low
+ 907.600000n V_low
+ 907.600001n V_low
+ 907.700000n V_low
+ 907.700001n V_low
+ 907.800000n V_low
+ 907.800001n V_low
+ 907.900000n V_low
+ 907.900001n V_low
+ 908.000000n V_low
+ 908.000001n V_low
+ 908.100000n V_low
+ 908.100001n V_low
+ 908.200000n V_low
+ 908.200001n V_low
+ 908.300000n V_low
+ 908.300001n V_low
+ 908.400000n V_low
+ 908.400001n V_low
+ 908.500000n V_low
+ 908.500001n V_low
+ 908.600000n V_low
+ 908.600001n V_low
+ 908.700000n V_low
+ 908.700001n V_low
+ 908.800000n V_low
+ 908.800001n V_low
+ 908.900000n V_low
+ 908.900001n V_low
+ 909.000000n V_low
+ 909.000001n V_hig
+ 909.100000n V_hig
+ 909.100001n V_hig
+ 909.200000n V_hig
+ 909.200001n V_hig
+ 909.300000n V_hig
+ 909.300001n V_hig
+ 909.400000n V_hig
+ 909.400001n V_hig
+ 909.500000n V_hig
+ 909.500001n V_hig
+ 909.600000n V_hig
+ 909.600001n V_hig
+ 909.700000n V_hig
+ 909.700001n V_hig
+ 909.800000n V_hig
+ 909.800001n V_hig
+ 909.900000n V_hig
+ 909.900001n V_hig
+ 910.000000n V_hig
+ 910.000001n V_hig
+ 910.100000n V_hig
+ 910.100001n V_hig
+ 910.200000n V_hig
+ 910.200001n V_hig
+ 910.300000n V_hig
+ 910.300001n V_hig
+ 910.400000n V_hig
+ 910.400001n V_hig
+ 910.500000n V_hig
+ 910.500001n V_hig
+ 910.600000n V_hig
+ 910.600001n V_hig
+ 910.700000n V_hig
+ 910.700001n V_hig
+ 910.800000n V_hig
+ 910.800001n V_hig
+ 910.900000n V_hig
+ 910.900001n V_hig
+ 911.000000n V_hig
+ 911.000001n V_hig
+ 911.100000n V_hig
+ 911.100001n V_hig
+ 911.200000n V_hig
+ 911.200001n V_hig
+ 911.300000n V_hig
+ 911.300001n V_hig
+ 911.400000n V_hig
+ 911.400001n V_hig
+ 911.500000n V_hig
+ 911.500001n V_hig
+ 911.600000n V_hig
+ 911.600001n V_hig
+ 911.700000n V_hig
+ 911.700001n V_hig
+ 911.800000n V_hig
+ 911.800001n V_hig
+ 911.900000n V_hig
+ 911.900001n V_hig
+ 912.000000n V_hig
+ 912.000001n V_hig
+ 912.100000n V_hig
+ 912.100001n V_hig
+ 912.200000n V_hig
+ 912.200001n V_hig
+ 912.300000n V_hig
+ 912.300001n V_hig
+ 912.400000n V_hig
+ 912.400001n V_hig
+ 912.500000n V_hig
+ 912.500001n V_hig
+ 912.600000n V_hig
+ 912.600001n V_hig
+ 912.700000n V_hig
+ 912.700001n V_hig
+ 912.800000n V_hig
+ 912.800001n V_hig
+ 912.900000n V_hig
+ 912.900001n V_hig
+ 913.000000n V_hig
+ 913.000001n V_hig
+ 913.100000n V_hig
+ 913.100001n V_hig
+ 913.200000n V_hig
+ 913.200001n V_hig
+ 913.300000n V_hig
+ 913.300001n V_hig
+ 913.400000n V_hig
+ 913.400001n V_hig
+ 913.500000n V_hig
+ 913.500001n V_hig
+ 913.600000n V_hig
+ 913.600001n V_hig
+ 913.700000n V_hig
+ 913.700001n V_hig
+ 913.800000n V_hig
+ 913.800001n V_hig
+ 913.900000n V_hig
+ 913.900001n V_hig
+ 914.000000n V_hig
+ 914.000001n V_hig
+ 914.100000n V_hig
+ 914.100001n V_hig
+ 914.200000n V_hig
+ 914.200001n V_hig
+ 914.300000n V_hig
+ 914.300001n V_hig
+ 914.400000n V_hig
+ 914.400001n V_hig
+ 914.500000n V_hig
+ 914.500001n V_hig
+ 914.600000n V_hig
+ 914.600001n V_hig
+ 914.700000n V_hig
+ 914.700001n V_hig
+ 914.800000n V_hig
+ 914.800001n V_hig
+ 914.900000n V_hig
+ 914.900001n V_hig
+ 915.000000n V_hig
+ 915.000001n V_hig
+ 915.100000n V_hig
+ 915.100001n V_hig
+ 915.200000n V_hig
+ 915.200001n V_hig
+ 915.300000n V_hig
+ 915.300001n V_hig
+ 915.400000n V_hig
+ 915.400001n V_hig
+ 915.500000n V_hig
+ 915.500001n V_hig
+ 915.600000n V_hig
+ 915.600001n V_hig
+ 915.700000n V_hig
+ 915.700001n V_hig
+ 915.800000n V_hig
+ 915.800001n V_hig
+ 915.900000n V_hig
+ 915.900001n V_hig
+ 916.000000n V_hig
+ 916.000001n V_hig
+ 916.100000n V_hig
+ 916.100001n V_hig
+ 916.200000n V_hig
+ 916.200001n V_hig
+ 916.300000n V_hig
+ 916.300001n V_hig
+ 916.400000n V_hig
+ 916.400001n V_hig
+ 916.500000n V_hig
+ 916.500001n V_hig
+ 916.600000n V_hig
+ 916.600001n V_hig
+ 916.700000n V_hig
+ 916.700001n V_hig
+ 916.800000n V_hig
+ 916.800001n V_hig
+ 916.900000n V_hig
+ 916.900001n V_hig
+ 917.000000n V_hig
+ 917.000001n V_low
+ 917.100000n V_low
+ 917.100001n V_low
+ 917.200000n V_low
+ 917.200001n V_low
+ 917.300000n V_low
+ 917.300001n V_low
+ 917.400000n V_low
+ 917.400001n V_low
+ 917.500000n V_low
+ 917.500001n V_low
+ 917.600000n V_low
+ 917.600001n V_low
+ 917.700000n V_low
+ 917.700001n V_low
+ 917.800000n V_low
+ 917.800001n V_low
+ 917.900000n V_low
+ 917.900001n V_low
+ 918.000000n V_low
+ 918.000001n V_hig
+ 918.100000n V_hig
+ 918.100001n V_hig
+ 918.200000n V_hig
+ 918.200001n V_hig
+ 918.300000n V_hig
+ 918.300001n V_hig
+ 918.400000n V_hig
+ 918.400001n V_hig
+ 918.500000n V_hig
+ 918.500001n V_hig
+ 918.600000n V_hig
+ 918.600001n V_hig
+ 918.700000n V_hig
+ 918.700001n V_hig
+ 918.800000n V_hig
+ 918.800001n V_hig
+ 918.900000n V_hig
+ 918.900001n V_hig
+ 919.000000n V_hig
+ 919.000001n V_hig
+ 919.100000n V_hig
+ 919.100001n V_hig
+ 919.200000n V_hig
+ 919.200001n V_hig
+ 919.300000n V_hig
+ 919.300001n V_hig
+ 919.400000n V_hig
+ 919.400001n V_hig
+ 919.500000n V_hig
+ 919.500001n V_hig
+ 919.600000n V_hig
+ 919.600001n V_hig
+ 919.700000n V_hig
+ 919.700001n V_hig
+ 919.800000n V_hig
+ 919.800001n V_hig
+ 919.900000n V_hig
+ 919.900001n V_hig
+ 920.000000n V_hig
+ 920.000001n V_hig
+ 920.100000n V_hig
+ 920.100001n V_hig
+ 920.200000n V_hig
+ 920.200001n V_hig
+ 920.300000n V_hig
+ 920.300001n V_hig
+ 920.400000n V_hig
+ 920.400001n V_hig
+ 920.500000n V_hig
+ 920.500001n V_hig
+ 920.600000n V_hig
+ 920.600001n V_hig
+ 920.700000n V_hig
+ 920.700001n V_hig
+ 920.800000n V_hig
+ 920.800001n V_hig
+ 920.900000n V_hig
+ 920.900001n V_hig
+ 921.000000n V_hig
+ 921.000001n V_low
+ 921.100000n V_low
+ 921.100001n V_low
+ 921.200000n V_low
+ 921.200001n V_low
+ 921.300000n V_low
+ 921.300001n V_low
+ 921.400000n V_low
+ 921.400001n V_low
+ 921.500000n V_low
+ 921.500001n V_low
+ 921.600000n V_low
+ 921.600001n V_low
+ 921.700000n V_low
+ 921.700001n V_low
+ 921.800000n V_low
+ 921.800001n V_low
+ 921.900000n V_low
+ 921.900001n V_low
+ 922.000000n V_low
+ 922.000001n V_low
+ 922.100000n V_low
+ 922.100001n V_low
+ 922.200000n V_low
+ 922.200001n V_low
+ 922.300000n V_low
+ 922.300001n V_low
+ 922.400000n V_low
+ 922.400001n V_low
+ 922.500000n V_low
+ 922.500001n V_low
+ 922.600000n V_low
+ 922.600001n V_low
+ 922.700000n V_low
+ 922.700001n V_low
+ 922.800000n V_low
+ 922.800001n V_low
+ 922.900000n V_low
+ 922.900001n V_low
+ 923.000000n V_low
+ 923.000001n V_hig
+ 923.100000n V_hig
+ 923.100001n V_hig
+ 923.200000n V_hig
+ 923.200001n V_hig
+ 923.300000n V_hig
+ 923.300001n V_hig
+ 923.400000n V_hig
+ 923.400001n V_hig
+ 923.500000n V_hig
+ 923.500001n V_hig
+ 923.600000n V_hig
+ 923.600001n V_hig
+ 923.700000n V_hig
+ 923.700001n V_hig
+ 923.800000n V_hig
+ 923.800001n V_hig
+ 923.900000n V_hig
+ 923.900001n V_hig
+ 924.000000n V_hig
+ 924.000001n V_hig
+ 924.100000n V_hig
+ 924.100001n V_hig
+ 924.200000n V_hig
+ 924.200001n V_hig
+ 924.300000n V_hig
+ 924.300001n V_hig
+ 924.400000n V_hig
+ 924.400001n V_hig
+ 924.500000n V_hig
+ 924.500001n V_hig
+ 924.600000n V_hig
+ 924.600001n V_hig
+ 924.700000n V_hig
+ 924.700001n V_hig
+ 924.800000n V_hig
+ 924.800001n V_hig
+ 924.900000n V_hig
+ 924.900001n V_hig
+ 925.000000n V_hig
+ 925.000001n V_low
+ 925.100000n V_low
+ 925.100001n V_low
+ 925.200000n V_low
+ 925.200001n V_low
+ 925.300000n V_low
+ 925.300001n V_low
+ 925.400000n V_low
+ 925.400001n V_low
+ 925.500000n V_low
+ 925.500001n V_low
+ 925.600000n V_low
+ 925.600001n V_low
+ 925.700000n V_low
+ 925.700001n V_low
+ 925.800000n V_low
+ 925.800001n V_low
+ 925.900000n V_low
+ 925.900001n V_low
+ 926.000000n V_low
+ 926.000001n V_low
+ 926.100000n V_low
+ 926.100001n V_low
+ 926.200000n V_low
+ 926.200001n V_low
+ 926.300000n V_low
+ 926.300001n V_low
+ 926.400000n V_low
+ 926.400001n V_low
+ 926.500000n V_low
+ 926.500001n V_low
+ 926.600000n V_low
+ 926.600001n V_low
+ 926.700000n V_low
+ 926.700001n V_low
+ 926.800000n V_low
+ 926.800001n V_low
+ 926.900000n V_low
+ 926.900001n V_low
+ 927.000000n V_low
+ 927.000001n V_low
+ 927.100000n V_low
+ 927.100001n V_low
+ 927.200000n V_low
+ 927.200001n V_low
+ 927.300000n V_low
+ 927.300001n V_low
+ 927.400000n V_low
+ 927.400001n V_low
+ 927.500000n V_low
+ 927.500001n V_low
+ 927.600000n V_low
+ 927.600001n V_low
+ 927.700000n V_low
+ 927.700001n V_low
+ 927.800000n V_low
+ 927.800001n V_low
+ 927.900000n V_low
+ 927.900001n V_low
+ 928.000000n V_low
+ 928.000001n V_hig
+ 928.100000n V_hig
+ 928.100001n V_hig
+ 928.200000n V_hig
+ 928.200001n V_hig
+ 928.300000n V_hig
+ 928.300001n V_hig
+ 928.400000n V_hig
+ 928.400001n V_hig
+ 928.500000n V_hig
+ 928.500001n V_hig
+ 928.600000n V_hig
+ 928.600001n V_hig
+ 928.700000n V_hig
+ 928.700001n V_hig
+ 928.800000n V_hig
+ 928.800001n V_hig
+ 928.900000n V_hig
+ 928.900001n V_hig
+ 929.000000n V_hig
+ 929.000001n V_low
+ 929.100000n V_low
+ 929.100001n V_low
+ 929.200000n V_low
+ 929.200001n V_low
+ 929.300000n V_low
+ 929.300001n V_low
+ 929.400000n V_low
+ 929.400001n V_low
+ 929.500000n V_low
+ 929.500001n V_low
+ 929.600000n V_low
+ 929.600001n V_low
+ 929.700000n V_low
+ 929.700001n V_low
+ 929.800000n V_low
+ 929.800001n V_low
+ 929.900000n V_low
+ 929.900001n V_low
+ 930.000000n V_low
+ 930.000001n V_hig
+ 930.100000n V_hig
+ 930.100001n V_hig
+ 930.200000n V_hig
+ 930.200001n V_hig
+ 930.300000n V_hig
+ 930.300001n V_hig
+ 930.400000n V_hig
+ 930.400001n V_hig
+ 930.500000n V_hig
+ 930.500001n V_hig
+ 930.600000n V_hig
+ 930.600001n V_hig
+ 930.700000n V_hig
+ 930.700001n V_hig
+ 930.800000n V_hig
+ 930.800001n V_hig
+ 930.900000n V_hig
+ 930.900001n V_hig
+ 931.000000n V_hig
+ 931.000001n V_hig
+ 931.100000n V_hig
+ 931.100001n V_hig
+ 931.200000n V_hig
+ 931.200001n V_hig
+ 931.300000n V_hig
+ 931.300001n V_hig
+ 931.400000n V_hig
+ 931.400001n V_hig
+ 931.500000n V_hig
+ 931.500001n V_hig
+ 931.600000n V_hig
+ 931.600001n V_hig
+ 931.700000n V_hig
+ 931.700001n V_hig
+ 931.800000n V_hig
+ 931.800001n V_hig
+ 931.900000n V_hig
+ 931.900001n V_hig
+ 932.000000n V_hig
+ 932.000001n V_low
+ 932.100000n V_low
+ 932.100001n V_low
+ 932.200000n V_low
+ 932.200001n V_low
+ 932.300000n V_low
+ 932.300001n V_low
+ 932.400000n V_low
+ 932.400001n V_low
+ 932.500000n V_low
+ 932.500001n V_low
+ 932.600000n V_low
+ 932.600001n V_low
+ 932.700000n V_low
+ 932.700001n V_low
+ 932.800000n V_low
+ 932.800001n V_low
+ 932.900000n V_low
+ 932.900001n V_low
+ 933.000000n V_low
+ 933.000001n V_low
+ 933.100000n V_low
+ 933.100001n V_low
+ 933.200000n V_low
+ 933.200001n V_low
+ 933.300000n V_low
+ 933.300001n V_low
+ 933.400000n V_low
+ 933.400001n V_low
+ 933.500000n V_low
+ 933.500001n V_low
+ 933.600000n V_low
+ 933.600001n V_low
+ 933.700000n V_low
+ 933.700001n V_low
+ 933.800000n V_low
+ 933.800001n V_low
+ 933.900000n V_low
+ 933.900001n V_low
+ 934.000000n V_low
+ 934.000001n V_low
+ 934.100000n V_low
+ 934.100001n V_low
+ 934.200000n V_low
+ 934.200001n V_low
+ 934.300000n V_low
+ 934.300001n V_low
+ 934.400000n V_low
+ 934.400001n V_low
+ 934.500000n V_low
+ 934.500001n V_low
+ 934.600000n V_low
+ 934.600001n V_low
+ 934.700000n V_low
+ 934.700001n V_low
+ 934.800000n V_low
+ 934.800001n V_low
+ 934.900000n V_low
+ 934.900001n V_low
+ 935.000000n V_low
+ 935.000001n V_hig
+ 935.100000n V_hig
+ 935.100001n V_hig
+ 935.200000n V_hig
+ 935.200001n V_hig
+ 935.300000n V_hig
+ 935.300001n V_hig
+ 935.400000n V_hig
+ 935.400001n V_hig
+ 935.500000n V_hig
+ 935.500001n V_hig
+ 935.600000n V_hig
+ 935.600001n V_hig
+ 935.700000n V_hig
+ 935.700001n V_hig
+ 935.800000n V_hig
+ 935.800001n V_hig
+ 935.900000n V_hig
+ 935.900001n V_hig
+ 936.000000n V_hig
+ 936.000001n V_low
+ 936.100000n V_low
+ 936.100001n V_low
+ 936.200000n V_low
+ 936.200001n V_low
+ 936.300000n V_low
+ 936.300001n V_low
+ 936.400000n V_low
+ 936.400001n V_low
+ 936.500000n V_low
+ 936.500001n V_low
+ 936.600000n V_low
+ 936.600001n V_low
+ 936.700000n V_low
+ 936.700001n V_low
+ 936.800000n V_low
+ 936.800001n V_low
+ 936.900000n V_low
+ 936.900001n V_low
+ 937.000000n V_low
+ 937.000001n V_hig
+ 937.100000n V_hig
+ 937.100001n V_hig
+ 937.200000n V_hig
+ 937.200001n V_hig
+ 937.300000n V_hig
+ 937.300001n V_hig
+ 937.400000n V_hig
+ 937.400001n V_hig
+ 937.500000n V_hig
+ 937.500001n V_hig
+ 937.600000n V_hig
+ 937.600001n V_hig
+ 937.700000n V_hig
+ 937.700001n V_hig
+ 937.800000n V_hig
+ 937.800001n V_hig
+ 937.900000n V_hig
+ 937.900001n V_hig
+ 938.000000n V_hig
+ 938.000001n V_low
+ 938.100000n V_low
+ 938.100001n V_low
+ 938.200000n V_low
+ 938.200001n V_low
+ 938.300000n V_low
+ 938.300001n V_low
+ 938.400000n V_low
+ 938.400001n V_low
+ 938.500000n V_low
+ 938.500001n V_low
+ 938.600000n V_low
+ 938.600001n V_low
+ 938.700000n V_low
+ 938.700001n V_low
+ 938.800000n V_low
+ 938.800001n V_low
+ 938.900000n V_low
+ 938.900001n V_low
+ 939.000000n V_low
+ 939.000001n V_low
+ 939.100000n V_low
+ 939.100001n V_low
+ 939.200000n V_low
+ 939.200001n V_low
+ 939.300000n V_low
+ 939.300001n V_low
+ 939.400000n V_low
+ 939.400001n V_low
+ 939.500000n V_low
+ 939.500001n V_low
+ 939.600000n V_low
+ 939.600001n V_low
+ 939.700000n V_low
+ 939.700001n V_low
+ 939.800000n V_low
+ 939.800001n V_low
+ 939.900000n V_low
+ 939.900001n V_low
+ 940.000000n V_low
+ 940.000001n V_low
+ 940.100000n V_low
+ 940.100001n V_low
+ 940.200000n V_low
+ 940.200001n V_low
+ 940.300000n V_low
+ 940.300001n V_low
+ 940.400000n V_low
+ 940.400001n V_low
+ 940.500000n V_low
+ 940.500001n V_low
+ 940.600000n V_low
+ 940.600001n V_low
+ 940.700000n V_low
+ 940.700001n V_low
+ 940.800000n V_low
+ 940.800001n V_low
+ 940.900000n V_low
+ 940.900001n V_low
+ 941.000000n V_low
+ 941.000001n V_hig
+ 941.100000n V_hig
+ 941.100001n V_hig
+ 941.200000n V_hig
+ 941.200001n V_hig
+ 941.300000n V_hig
+ 941.300001n V_hig
+ 941.400000n V_hig
+ 941.400001n V_hig
+ 941.500000n V_hig
+ 941.500001n V_hig
+ 941.600000n V_hig
+ 941.600001n V_hig
+ 941.700000n V_hig
+ 941.700001n V_hig
+ 941.800000n V_hig
+ 941.800001n V_hig
+ 941.900000n V_hig
+ 941.900001n V_hig
+ 942.000000n V_hig
+ 942.000001n V_low
+ 942.100000n V_low
+ 942.100001n V_low
+ 942.200000n V_low
+ 942.200001n V_low
+ 942.300000n V_low
+ 942.300001n V_low
+ 942.400000n V_low
+ 942.400001n V_low
+ 942.500000n V_low
+ 942.500001n V_low
+ 942.600000n V_low
+ 942.600001n V_low
+ 942.700000n V_low
+ 942.700001n V_low
+ 942.800000n V_low
+ 942.800001n V_low
+ 942.900000n V_low
+ 942.900001n V_low
+ 943.000000n V_low
+ 943.000001n V_low
+ 943.100000n V_low
+ 943.100001n V_low
+ 943.200000n V_low
+ 943.200001n V_low
+ 943.300000n V_low
+ 943.300001n V_low
+ 943.400000n V_low
+ 943.400001n V_low
+ 943.500000n V_low
+ 943.500001n V_low
+ 943.600000n V_low
+ 943.600001n V_low
+ 943.700000n V_low
+ 943.700001n V_low
+ 943.800000n V_low
+ 943.800001n V_low
+ 943.900000n V_low
+ 943.900001n V_low
+ 944.000000n V_low
+ 944.000001n V_hig
+ 944.100000n V_hig
+ 944.100001n V_hig
+ 944.200000n V_hig
+ 944.200001n V_hig
+ 944.300000n V_hig
+ 944.300001n V_hig
+ 944.400000n V_hig
+ 944.400001n V_hig
+ 944.500000n V_hig
+ 944.500001n V_hig
+ 944.600000n V_hig
+ 944.600001n V_hig
+ 944.700000n V_hig
+ 944.700001n V_hig
+ 944.800000n V_hig
+ 944.800001n V_hig
+ 944.900000n V_hig
+ 944.900001n V_hig
+ 945.000000n V_hig
+ 945.000001n V_hig
+ 945.100000n V_hig
+ 945.100001n V_hig
+ 945.200000n V_hig
+ 945.200001n V_hig
+ 945.300000n V_hig
+ 945.300001n V_hig
+ 945.400000n V_hig
+ 945.400001n V_hig
+ 945.500000n V_hig
+ 945.500001n V_hig
+ 945.600000n V_hig
+ 945.600001n V_hig
+ 945.700000n V_hig
+ 945.700001n V_hig
+ 945.800000n V_hig
+ 945.800001n V_hig
+ 945.900000n V_hig
+ 945.900001n V_hig
+ 946.000000n V_hig
+ 946.000001n V_low
+ 946.100000n V_low
+ 946.100001n V_low
+ 946.200000n V_low
+ 946.200001n V_low
+ 946.300000n V_low
+ 946.300001n V_low
+ 946.400000n V_low
+ 946.400001n V_low
+ 946.500000n V_low
+ 946.500001n V_low
+ 946.600000n V_low
+ 946.600001n V_low
+ 946.700000n V_low
+ 946.700001n V_low
+ 946.800000n V_low
+ 946.800001n V_low
+ 946.900000n V_low
+ 946.900001n V_low
+ 947.000000n V_low
+ 947.000001n V_hig
+ 947.100000n V_hig
+ 947.100001n V_hig
+ 947.200000n V_hig
+ 947.200001n V_hig
+ 947.300000n V_hig
+ 947.300001n V_hig
+ 947.400000n V_hig
+ 947.400001n V_hig
+ 947.500000n V_hig
+ 947.500001n V_hig
+ 947.600000n V_hig
+ 947.600001n V_hig
+ 947.700000n V_hig
+ 947.700001n V_hig
+ 947.800000n V_hig
+ 947.800001n V_hig
+ 947.900000n V_hig
+ 947.900001n V_hig
+ 948.000000n V_hig
+ 948.000001n V_low
+ 948.100000n V_low
+ 948.100001n V_low
+ 948.200000n V_low
+ 948.200001n V_low
+ 948.300000n V_low
+ 948.300001n V_low
+ 948.400000n V_low
+ 948.400001n V_low
+ 948.500000n V_low
+ 948.500001n V_low
+ 948.600000n V_low
+ 948.600001n V_low
+ 948.700000n V_low
+ 948.700001n V_low
+ 948.800000n V_low
+ 948.800001n V_low
+ 948.900000n V_low
+ 948.900001n V_low
+ 949.000000n V_low
+ 949.000001n V_low
+ 949.100000n V_low
+ 949.100001n V_low
+ 949.200000n V_low
+ 949.200001n V_low
+ 949.300000n V_low
+ 949.300001n V_low
+ 949.400000n V_low
+ 949.400001n V_low
+ 949.500000n V_low
+ 949.500001n V_low
+ 949.600000n V_low
+ 949.600001n V_low
+ 949.700000n V_low
+ 949.700001n V_low
+ 949.800000n V_low
+ 949.800001n V_low
+ 949.900000n V_low
+ 949.900001n V_low
+ 950.000000n V_low
+ 950.000001n V_hig
+ 950.100000n V_hig
+ 950.100001n V_hig
+ 950.200000n V_hig
+ 950.200001n V_hig
+ 950.300000n V_hig
+ 950.300001n V_hig
+ 950.400000n V_hig
+ 950.400001n V_hig
+ 950.500000n V_hig
+ 950.500001n V_hig
+ 950.600000n V_hig
+ 950.600001n V_hig
+ 950.700000n V_hig
+ 950.700001n V_hig
+ 950.800000n V_hig
+ 950.800001n V_hig
+ 950.900000n V_hig
+ 950.900001n V_hig
+ 951.000000n V_hig
+ 951.000001n V_low
+ 951.100000n V_low
+ 951.100001n V_low
+ 951.200000n V_low
+ 951.200001n V_low
+ 951.300000n V_low
+ 951.300001n V_low
+ 951.400000n V_low
+ 951.400001n V_low
+ 951.500000n V_low
+ 951.500001n V_low
+ 951.600000n V_low
+ 951.600001n V_low
+ 951.700000n V_low
+ 951.700001n V_low
+ 951.800000n V_low
+ 951.800001n V_low
+ 951.900000n V_low
+ 951.900001n V_low
+ 952.000000n V_low
+ 952.000001n V_low
+ 952.100000n V_low
+ 952.100001n V_low
+ 952.200000n V_low
+ 952.200001n V_low
+ 952.300000n V_low
+ 952.300001n V_low
+ 952.400000n V_low
+ 952.400001n V_low
+ 952.500000n V_low
+ 952.500001n V_low
+ 952.600000n V_low
+ 952.600001n V_low
+ 952.700000n V_low
+ 952.700001n V_low
+ 952.800000n V_low
+ 952.800001n V_low
+ 952.900000n V_low
+ 952.900001n V_low
+ 953.000000n V_low
+ 953.000001n V_hig
+ 953.100000n V_hig
+ 953.100001n V_hig
+ 953.200000n V_hig
+ 953.200001n V_hig
+ 953.300000n V_hig
+ 953.300001n V_hig
+ 953.400000n V_hig
+ 953.400001n V_hig
+ 953.500000n V_hig
+ 953.500001n V_hig
+ 953.600000n V_hig
+ 953.600001n V_hig
+ 953.700000n V_hig
+ 953.700001n V_hig
+ 953.800000n V_hig
+ 953.800001n V_hig
+ 953.900000n V_hig
+ 953.900001n V_hig
+ 954.000000n V_hig
+ 954.000001n V_low
+ 954.100000n V_low
+ 954.100001n V_low
+ 954.200000n V_low
+ 954.200001n V_low
+ 954.300000n V_low
+ 954.300001n V_low
+ 954.400000n V_low
+ 954.400001n V_low
+ 954.500000n V_low
+ 954.500001n V_low
+ 954.600000n V_low
+ 954.600001n V_low
+ 954.700000n V_low
+ 954.700001n V_low
+ 954.800000n V_low
+ 954.800001n V_low
+ 954.900000n V_low
+ 954.900001n V_low
+ 955.000000n V_low
+ 955.000001n V_hig
+ 955.100000n V_hig
+ 955.100001n V_hig
+ 955.200000n V_hig
+ 955.200001n V_hig
+ 955.300000n V_hig
+ 955.300001n V_hig
+ 955.400000n V_hig
+ 955.400001n V_hig
+ 955.500000n V_hig
+ 955.500001n V_hig
+ 955.600000n V_hig
+ 955.600001n V_hig
+ 955.700000n V_hig
+ 955.700001n V_hig
+ 955.800000n V_hig
+ 955.800001n V_hig
+ 955.900000n V_hig
+ 955.900001n V_hig
+ 956.000000n V_hig
+ 956.000001n V_low
+ 956.100000n V_low
+ 956.100001n V_low
+ 956.200000n V_low
+ 956.200001n V_low
+ 956.300000n V_low
+ 956.300001n V_low
+ 956.400000n V_low
+ 956.400001n V_low
+ 956.500000n V_low
+ 956.500001n V_low
+ 956.600000n V_low
+ 956.600001n V_low
+ 956.700000n V_low
+ 956.700001n V_low
+ 956.800000n V_low
+ 956.800001n V_low
+ 956.900000n V_low
+ 956.900001n V_low
+ 957.000000n V_low
+ 957.000001n V_hig
+ 957.100000n V_hig
+ 957.100001n V_hig
+ 957.200000n V_hig
+ 957.200001n V_hig
+ 957.300000n V_hig
+ 957.300001n V_hig
+ 957.400000n V_hig
+ 957.400001n V_hig
+ 957.500000n V_hig
+ 957.500001n V_hig
+ 957.600000n V_hig
+ 957.600001n V_hig
+ 957.700000n V_hig
+ 957.700001n V_hig
+ 957.800000n V_hig
+ 957.800001n V_hig
+ 957.900000n V_hig
+ 957.900001n V_hig
+ 958.000000n V_hig
+ 958.000001n V_low
+ 958.100000n V_low
+ 958.100001n V_low
+ 958.200000n V_low
+ 958.200001n V_low
+ 958.300000n V_low
+ 958.300001n V_low
+ 958.400000n V_low
+ 958.400001n V_low
+ 958.500000n V_low
+ 958.500001n V_low
+ 958.600000n V_low
+ 958.600001n V_low
+ 958.700000n V_low
+ 958.700001n V_low
+ 958.800000n V_low
+ 958.800001n V_low
+ 958.900000n V_low
+ 958.900001n V_low
+ 959.000000n V_low
+ 959.000001n V_low
+ 959.100000n V_low
+ 959.100001n V_low
+ 959.200000n V_low
+ 959.200001n V_low
+ 959.300000n V_low
+ 959.300001n V_low
+ 959.400000n V_low
+ 959.400001n V_low
+ 959.500000n V_low
+ 959.500001n V_low
+ 959.600000n V_low
+ 959.600001n V_low
+ 959.700000n V_low
+ 959.700001n V_low
+ 959.800000n V_low
+ 959.800001n V_low
+ 959.900000n V_low
+ 959.900001n V_low
+ 960.000000n V_low
+ 960.000001n V_hig
+ 960.100000n V_hig
+ 960.100001n V_hig
+ 960.200000n V_hig
+ 960.200001n V_hig
+ 960.300000n V_hig
+ 960.300001n V_hig
+ 960.400000n V_hig
+ 960.400001n V_hig
+ 960.500000n V_hig
+ 960.500001n V_hig
+ 960.600000n V_hig
+ 960.600001n V_hig
+ 960.700000n V_hig
+ 960.700001n V_hig
+ 960.800000n V_hig
+ 960.800001n V_hig
+ 960.900000n V_hig
+ 960.900001n V_hig
+ 961.000000n V_hig
+ 961.000001n V_hig
+ 961.100000n V_hig
+ 961.100001n V_hig
+ 961.200000n V_hig
+ 961.200001n V_hig
+ 961.300000n V_hig
+ 961.300001n V_hig
+ 961.400000n V_hig
+ 961.400001n V_hig
+ 961.500000n V_hig
+ 961.500001n V_hig
+ 961.600000n V_hig
+ 961.600001n V_hig
+ 961.700000n V_hig
+ 961.700001n V_hig
+ 961.800000n V_hig
+ 961.800001n V_hig
+ 961.900000n V_hig
+ 961.900001n V_hig
+ 962.000000n V_hig
+ 962.000001n V_low
+ 962.100000n V_low
+ 962.100001n V_low
+ 962.200000n V_low
+ 962.200001n V_low
+ 962.300000n V_low
+ 962.300001n V_low
+ 962.400000n V_low
+ 962.400001n V_low
+ 962.500000n V_low
+ 962.500001n V_low
+ 962.600000n V_low
+ 962.600001n V_low
+ 962.700000n V_low
+ 962.700001n V_low
+ 962.800000n V_low
+ 962.800001n V_low
+ 962.900000n V_low
+ 962.900001n V_low
+ 963.000000n V_low
+ 963.000001n V_low
+ 963.100000n V_low
+ 963.100001n V_low
+ 963.200000n V_low
+ 963.200001n V_low
+ 963.300000n V_low
+ 963.300001n V_low
+ 963.400000n V_low
+ 963.400001n V_low
+ 963.500000n V_low
+ 963.500001n V_low
+ 963.600000n V_low
+ 963.600001n V_low
+ 963.700000n V_low
+ 963.700001n V_low
+ 963.800000n V_low
+ 963.800001n V_low
+ 963.900000n V_low
+ 963.900001n V_low
+ 964.000000n V_low
+ 964.000001n V_low
+ 964.100000n V_low
+ 964.100001n V_low
+ 964.200000n V_low
+ 964.200001n V_low
+ 964.300000n V_low
+ 964.300001n V_low
+ 964.400000n V_low
+ 964.400001n V_low
+ 964.500000n V_low
+ 964.500001n V_low
+ 964.600000n V_low
+ 964.600001n V_low
+ 964.700000n V_low
+ 964.700001n V_low
+ 964.800000n V_low
+ 964.800001n V_low
+ 964.900000n V_low
+ 964.900001n V_low
+ 965.000000n V_low
+ 965.000001n V_hig
+ 965.100000n V_hig
+ 965.100001n V_hig
+ 965.200000n V_hig
+ 965.200001n V_hig
+ 965.300000n V_hig
+ 965.300001n V_hig
+ 965.400000n V_hig
+ 965.400001n V_hig
+ 965.500000n V_hig
+ 965.500001n V_hig
+ 965.600000n V_hig
+ 965.600001n V_hig
+ 965.700000n V_hig
+ 965.700001n V_hig
+ 965.800000n V_hig
+ 965.800001n V_hig
+ 965.900000n V_hig
+ 965.900001n V_hig
+ 966.000000n V_hig
+ 966.000001n V_low
+ 966.100000n V_low
+ 966.100001n V_low
+ 966.200000n V_low
+ 966.200001n V_low
+ 966.300000n V_low
+ 966.300001n V_low
+ 966.400000n V_low
+ 966.400001n V_low
+ 966.500000n V_low
+ 966.500001n V_low
+ 966.600000n V_low
+ 966.600001n V_low
+ 966.700000n V_low
+ 966.700001n V_low
+ 966.800000n V_low
+ 966.800001n V_low
+ 966.900000n V_low
+ 966.900001n V_low
+ 967.000000n V_low
+ 967.000001n V_hig
+ 967.100000n V_hig
+ 967.100001n V_hig
+ 967.200000n V_hig
+ 967.200001n V_hig
+ 967.300000n V_hig
+ 967.300001n V_hig
+ 967.400000n V_hig
+ 967.400001n V_hig
+ 967.500000n V_hig
+ 967.500001n V_hig
+ 967.600000n V_hig
+ 967.600001n V_hig
+ 967.700000n V_hig
+ 967.700001n V_hig
+ 967.800000n V_hig
+ 967.800001n V_hig
+ 967.900000n V_hig
+ 967.900001n V_hig
+ 968.000000n V_hig
+ 968.000001n V_hig
+ 968.100000n V_hig
+ 968.100001n V_hig
+ 968.200000n V_hig
+ 968.200001n V_hig
+ 968.300000n V_hig
+ 968.300001n V_hig
+ 968.400000n V_hig
+ 968.400001n V_hig
+ 968.500000n V_hig
+ 968.500001n V_hig
+ 968.600000n V_hig
+ 968.600001n V_hig
+ 968.700000n V_hig
+ 968.700001n V_hig
+ 968.800000n V_hig
+ 968.800001n V_hig
+ 968.900000n V_hig
+ 968.900001n V_hig
+ 969.000000n V_hig
+ 969.000001n V_low
+ 969.100000n V_low
+ 969.100001n V_low
+ 969.200000n V_low
+ 969.200001n V_low
+ 969.300000n V_low
+ 969.300001n V_low
+ 969.400000n V_low
+ 969.400001n V_low
+ 969.500000n V_low
+ 969.500001n V_low
+ 969.600000n V_low
+ 969.600001n V_low
+ 969.700000n V_low
+ 969.700001n V_low
+ 969.800000n V_low
+ 969.800001n V_low
+ 969.900000n V_low
+ 969.900001n V_low
+ 970.000000n V_low
+ 970.000001n V_hig
+ 970.100000n V_hig
+ 970.100001n V_hig
+ 970.200000n V_hig
+ 970.200001n V_hig
+ 970.300000n V_hig
+ 970.300001n V_hig
+ 970.400000n V_hig
+ 970.400001n V_hig
+ 970.500000n V_hig
+ 970.500001n V_hig
+ 970.600000n V_hig
+ 970.600001n V_hig
+ 970.700000n V_hig
+ 970.700001n V_hig
+ 970.800000n V_hig
+ 970.800001n V_hig
+ 970.900000n V_hig
+ 970.900001n V_hig
+ 971.000000n V_hig
+ 971.000001n V_hig
+ 971.100000n V_hig
+ 971.100001n V_hig
+ 971.200000n V_hig
+ 971.200001n V_hig
+ 971.300000n V_hig
+ 971.300001n V_hig
+ 971.400000n V_hig
+ 971.400001n V_hig
+ 971.500000n V_hig
+ 971.500001n V_hig
+ 971.600000n V_hig
+ 971.600001n V_hig
+ 971.700000n V_hig
+ 971.700001n V_hig
+ 971.800000n V_hig
+ 971.800001n V_hig
+ 971.900000n V_hig
+ 971.900001n V_hig
+ 972.000000n V_hig
+ 972.000001n V_low
+ 972.100000n V_low
+ 972.100001n V_low
+ 972.200000n V_low
+ 972.200001n V_low
+ 972.300000n V_low
+ 972.300001n V_low
+ 972.400000n V_low
+ 972.400001n V_low
+ 972.500000n V_low
+ 972.500001n V_low
+ 972.600000n V_low
+ 972.600001n V_low
+ 972.700000n V_low
+ 972.700001n V_low
+ 972.800000n V_low
+ 972.800001n V_low
+ 972.900000n V_low
+ 972.900001n V_low
+ 973.000000n V_low
+ 973.000001n V_hig
+ 973.100000n V_hig
+ 973.100001n V_hig
+ 973.200000n V_hig
+ 973.200001n V_hig
+ 973.300000n V_hig
+ 973.300001n V_hig
+ 973.400000n V_hig
+ 973.400001n V_hig
+ 973.500000n V_hig
+ 973.500001n V_hig
+ 973.600000n V_hig
+ 973.600001n V_hig
+ 973.700000n V_hig
+ 973.700001n V_hig
+ 973.800000n V_hig
+ 973.800001n V_hig
+ 973.900000n V_hig
+ 973.900001n V_hig
+ 974.000000n V_hig
+ 974.000001n V_low
+ 974.100000n V_low
+ 974.100001n V_low
+ 974.200000n V_low
+ 974.200001n V_low
+ 974.300000n V_low
+ 974.300001n V_low
+ 974.400000n V_low
+ 974.400001n V_low
+ 974.500000n V_low
+ 974.500001n V_low
+ 974.600000n V_low
+ 974.600001n V_low
+ 974.700000n V_low
+ 974.700001n V_low
+ 974.800000n V_low
+ 974.800001n V_low
+ 974.900000n V_low
+ 974.900001n V_low
+ 975.000000n V_low
+ 975.000001n V_hig
+ 975.100000n V_hig
+ 975.100001n V_hig
+ 975.200000n V_hig
+ 975.200001n V_hig
+ 975.300000n V_hig
+ 975.300001n V_hig
+ 975.400000n V_hig
+ 975.400001n V_hig
+ 975.500000n V_hig
+ 975.500001n V_hig
+ 975.600000n V_hig
+ 975.600001n V_hig
+ 975.700000n V_hig
+ 975.700001n V_hig
+ 975.800000n V_hig
+ 975.800001n V_hig
+ 975.900000n V_hig
+ 975.900001n V_hig
+ 976.000000n V_hig
+ 976.000001n V_hig
+ 976.100000n V_hig
+ 976.100001n V_hig
+ 976.200000n V_hig
+ 976.200001n V_hig
+ 976.300000n V_hig
+ 976.300001n V_hig
+ 976.400000n V_hig
+ 976.400001n V_hig
+ 976.500000n V_hig
+ 976.500001n V_hig
+ 976.600000n V_hig
+ 976.600001n V_hig
+ 976.700000n V_hig
+ 976.700001n V_hig
+ 976.800000n V_hig
+ 976.800001n V_hig
+ 976.900000n V_hig
+ 976.900001n V_hig
+ 977.000000n V_hig
+ 977.000001n V_low
+ 977.100000n V_low
+ 977.100001n V_low
+ 977.200000n V_low
+ 977.200001n V_low
+ 977.300000n V_low
+ 977.300001n V_low
+ 977.400000n V_low
+ 977.400001n V_low
+ 977.500000n V_low
+ 977.500001n V_low
+ 977.600000n V_low
+ 977.600001n V_low
+ 977.700000n V_low
+ 977.700001n V_low
+ 977.800000n V_low
+ 977.800001n V_low
+ 977.900000n V_low
+ 977.900001n V_low
+ 978.000000n V_low
+ 978.000001n V_low
+ 978.100000n V_low
+ 978.100001n V_low
+ 978.200000n V_low
+ 978.200001n V_low
+ 978.300000n V_low
+ 978.300001n V_low
+ 978.400000n V_low
+ 978.400001n V_low
+ 978.500000n V_low
+ 978.500001n V_low
+ 978.600000n V_low
+ 978.600001n V_low
+ 978.700000n V_low
+ 978.700001n V_low
+ 978.800000n V_low
+ 978.800001n V_low
+ 978.900000n V_low
+ 978.900001n V_low
+ 979.000000n V_low
+ 979.000001n V_low
+ 979.100000n V_low
+ 979.100001n V_low
+ 979.200000n V_low
+ 979.200001n V_low
+ 979.300000n V_low
+ 979.300001n V_low
+ 979.400000n V_low
+ 979.400001n V_low
+ 979.500000n V_low
+ 979.500001n V_low
+ 979.600000n V_low
+ 979.600001n V_low
+ 979.700000n V_low
+ 979.700001n V_low
+ 979.800000n V_low
+ 979.800001n V_low
+ 979.900000n V_low
+ 979.900001n V_low
+ 980.000000n V_low
+ 980.000001n V_hig
+ 980.100000n V_hig
+ 980.100001n V_hig
+ 980.200000n V_hig
+ 980.200001n V_hig
+ 980.300000n V_hig
+ 980.300001n V_hig
+ 980.400000n V_hig
+ 980.400001n V_hig
+ 980.500000n V_hig
+ 980.500001n V_hig
+ 980.600000n V_hig
+ 980.600001n V_hig
+ 980.700000n V_hig
+ 980.700001n V_hig
+ 980.800000n V_hig
+ 980.800001n V_hig
+ 980.900000n V_hig
+ 980.900001n V_hig
+ 981.000000n V_hig
+ 981.000001n V_hig
+ 981.100000n V_hig
+ 981.100001n V_hig
+ 981.200000n V_hig
+ 981.200001n V_hig
+ 981.300000n V_hig
+ 981.300001n V_hig
+ 981.400000n V_hig
+ 981.400001n V_hig
+ 981.500000n V_hig
+ 981.500001n V_hig
+ 981.600000n V_hig
+ 981.600001n V_hig
+ 981.700000n V_hig
+ 981.700001n V_hig
+ 981.800000n V_hig
+ 981.800001n V_hig
+ 981.900000n V_hig
+ 981.900001n V_hig
+ 982.000000n V_hig
+ 982.000001n V_hig
+ 982.100000n V_hig
+ 982.100001n V_hig
+ 982.200000n V_hig
+ 982.200001n V_hig
+ 982.300000n V_hig
+ 982.300001n V_hig
+ 982.400000n V_hig
+ 982.400001n V_hig
+ 982.500000n V_hig
+ 982.500001n V_hig
+ 982.600000n V_hig
+ 982.600001n V_hig
+ 982.700000n V_hig
+ 982.700001n V_hig
+ 982.800000n V_hig
+ 982.800001n V_hig
+ 982.900000n V_hig
+ 982.900001n V_hig
+ 983.000000n V_hig
+ 983.000001n V_hig
+ 983.100000n V_hig
+ 983.100001n V_hig
+ 983.200000n V_hig
+ 983.200001n V_hig
+ 983.300000n V_hig
+ 983.300001n V_hig
+ 983.400000n V_hig
+ 983.400001n V_hig
+ 983.500000n V_hig
+ 983.500001n V_hig
+ 983.600000n V_hig
+ 983.600001n V_hig
+ 983.700000n V_hig
+ 983.700001n V_hig
+ 983.800000n V_hig
+ 983.800001n V_hig
+ 983.900000n V_hig
+ 983.900001n V_hig
+ 984.000000n V_hig
+ 984.000001n V_hig
+ 984.100000n V_hig
+ 984.100001n V_hig
+ 984.200000n V_hig
+ 984.200001n V_hig
+ 984.300000n V_hig
+ 984.300001n V_hig
+ 984.400000n V_hig
+ 984.400001n V_hig
+ 984.500000n V_hig
+ 984.500001n V_hig
+ 984.600000n V_hig
+ 984.600001n V_hig
+ 984.700000n V_hig
+ 984.700001n V_hig
+ 984.800000n V_hig
+ 984.800001n V_hig
+ 984.900000n V_hig
+ 984.900001n V_hig
+ 985.000000n V_hig
+ 985.000001n V_hig
+ 985.100000n V_hig
+ 985.100001n V_hig
+ 985.200000n V_hig
+ 985.200001n V_hig
+ 985.300000n V_hig
+ 985.300001n V_hig
+ 985.400000n V_hig
+ 985.400001n V_hig
+ 985.500000n V_hig
+ 985.500001n V_hig
+ 985.600000n V_hig
+ 985.600001n V_hig
+ 985.700000n V_hig
+ 985.700001n V_hig
+ 985.800000n V_hig
+ 985.800001n V_hig
+ 985.900000n V_hig
+ 985.900001n V_hig
+ 986.000000n V_hig
+ 986.000001n V_hig
+ 986.100000n V_hig
+ 986.100001n V_hig
+ 986.200000n V_hig
+ 986.200001n V_hig
+ 986.300000n V_hig
+ 986.300001n V_hig
+ 986.400000n V_hig
+ 986.400001n V_hig
+ 986.500000n V_hig
+ 986.500001n V_hig
+ 986.600000n V_hig
+ 986.600001n V_hig
+ 986.700000n V_hig
+ 986.700001n V_hig
+ 986.800000n V_hig
+ 986.800001n V_hig
+ 986.900000n V_hig
+ 986.900001n V_hig
+ 987.000000n V_hig
+ 987.000001n V_hig
+ 987.100000n V_hig
+ 987.100001n V_hig
+ 987.200000n V_hig
+ 987.200001n V_hig
+ 987.300000n V_hig
+ 987.300001n V_hig
+ 987.400000n V_hig
+ 987.400001n V_hig
+ 987.500000n V_hig
+ 987.500001n V_hig
+ 987.600000n V_hig
+ 987.600001n V_hig
+ 987.700000n V_hig
+ 987.700001n V_hig
+ 987.800000n V_hig
+ 987.800001n V_hig
+ 987.900000n V_hig
+ 987.900001n V_hig
+ 988.000000n V_hig
+ 988.000001n V_hig
+ 988.100000n V_hig
+ 988.100001n V_hig
+ 988.200000n V_hig
+ 988.200001n V_hig
+ 988.300000n V_hig
+ 988.300001n V_hig
+ 988.400000n V_hig
+ 988.400001n V_hig
+ 988.500000n V_hig
+ 988.500001n V_hig
+ 988.600000n V_hig
+ 988.600001n V_hig
+ 988.700000n V_hig
+ 988.700001n V_hig
+ 988.800000n V_hig
+ 988.800001n V_hig
+ 988.900000n V_hig
+ 988.900001n V_hig
+ 989.000000n V_hig
+ 989.000001n V_hig
+ 989.100000n V_hig
+ 989.100001n V_hig
+ 989.200000n V_hig
+ 989.200001n V_hig
+ 989.300000n V_hig
+ 989.300001n V_hig
+ 989.400000n V_hig
+ 989.400001n V_hig
+ 989.500000n V_hig
+ 989.500001n V_hig
+ 989.600000n V_hig
+ 989.600001n V_hig
+ 989.700000n V_hig
+ 989.700001n V_hig
+ 989.800000n V_hig
+ 989.800001n V_hig
+ 989.900000n V_hig
+ 989.900001n V_hig
+ 990.000000n V_hig
+ 990.000001n V_low
+ 990.100000n V_low
+ 990.100001n V_low
+ 990.200000n V_low
+ 990.200001n V_low
+ 990.300000n V_low
+ 990.300001n V_low
+ 990.400000n V_low
+ 990.400001n V_low
+ 990.500000n V_low
+ 990.500001n V_low
+ 990.600000n V_low
+ 990.600001n V_low
+ 990.700000n V_low
+ 990.700001n V_low
+ 990.800000n V_low
+ 990.800001n V_low
+ 990.900000n V_low
+ 990.900001n V_low
+ 991.000000n V_low
+ 991.000001n V_hig
+ 991.100000n V_hig
+ 991.100001n V_hig
+ 991.200000n V_hig
+ 991.200001n V_hig
+ 991.300000n V_hig
+ 991.300001n V_hig
+ 991.400000n V_hig
+ 991.400001n V_hig
+ 991.500000n V_hig
+ 991.500001n V_hig
+ 991.600000n V_hig
+ 991.600001n V_hig
+ 991.700000n V_hig
+ 991.700001n V_hig
+ 991.800000n V_hig
+ 991.800001n V_hig
+ 991.900000n V_hig
+ 991.900001n V_hig
+ 992.000000n V_hig
+ 992.000001n V_hig
+ 992.100000n V_hig
+ 992.100001n V_hig
+ 992.200000n V_hig
+ 992.200001n V_hig
+ 992.300000n V_hig
+ 992.300001n V_hig
+ 992.400000n V_hig
+ 992.400001n V_hig
+ 992.500000n V_hig
+ 992.500001n V_hig
+ 992.600000n V_hig
+ 992.600001n V_hig
+ 992.700000n V_hig
+ 992.700001n V_hig
+ 992.800000n V_hig
+ 992.800001n V_hig
+ 992.900000n V_hig
+ 992.900001n V_hig
+ 993.000000n V_hig
+ 993.000001n V_hig
+ 993.100000n V_hig
+ 993.100001n V_hig
+ 993.200000n V_hig
+ 993.200001n V_hig
+ 993.300000n V_hig
+ 993.300001n V_hig
+ 993.400000n V_hig
+ 993.400001n V_hig
+ 993.500000n V_hig
+ 993.500001n V_hig
+ 993.600000n V_hig
+ 993.600001n V_hig
+ 993.700000n V_hig
+ 993.700001n V_hig
+ 993.800000n V_hig
+ 993.800001n V_hig
+ 993.900000n V_hig
+ 993.900001n V_hig
+ 994.000000n V_hig
+ 994.000001n V_hig
+ 994.100000n V_hig
+ 994.100001n V_hig
+ 994.200000n V_hig
+ 994.200001n V_hig
+ 994.300000n V_hig
+ 994.300001n V_hig
+ 994.400000n V_hig
+ 994.400001n V_hig
+ 994.500000n V_hig
+ 994.500001n V_hig
+ 994.600000n V_hig
+ 994.600001n V_hig
+ 994.700000n V_hig
+ 994.700001n V_hig
+ 994.800000n V_hig
+ 994.800001n V_hig
+ 994.900000n V_hig
+ 994.900001n V_hig
+ 995.000000n V_hig
+ 995.000001n V_low
+ 995.100000n V_low
+ 995.100001n V_low
+ 995.200000n V_low
+ 995.200001n V_low
+ 995.300000n V_low
+ 995.300001n V_low
+ 995.400000n V_low
+ 995.400001n V_low
+ 995.500000n V_low
+ 995.500001n V_low
+ 995.600000n V_low
+ 995.600001n V_low
+ 995.700000n V_low
+ 995.700001n V_low
+ 995.800000n V_low
+ 995.800001n V_low
+ 995.900000n V_low
+ 995.900001n V_low
+ 996.000000n V_low
+ 996.000001n V_hig
+ 996.100000n V_hig
+ 996.100001n V_hig
+ 996.200000n V_hig
+ 996.200001n V_hig
+ 996.300000n V_hig
+ 996.300001n V_hig
+ 996.400000n V_hig
+ 996.400001n V_hig
+ 996.500000n V_hig
+ 996.500001n V_hig
+ 996.600000n V_hig
+ 996.600001n V_hig
+ 996.700000n V_hig
+ 996.700001n V_hig
+ 996.800000n V_hig
+ 996.800001n V_hig
+ 996.900000n V_hig
+ 996.900001n V_hig
+ 997.000000n V_hig
+ 997.000001n V_low
+ 997.100000n V_low
+ 997.100001n V_low
+ 997.200000n V_low
+ 997.200001n V_low
+ 997.300000n V_low
+ 997.300001n V_low
+ 997.400000n V_low
+ 997.400001n V_low
+ 997.500000n V_low
+ 997.500001n V_low
+ 997.600000n V_low
+ 997.600001n V_low
+ 997.700000n V_low
+ 997.700001n V_low
+ 997.800000n V_low
+ 997.800001n V_low
+ 997.900000n V_low
+ 997.900001n V_low
+ 998.000000n V_low
+ 998.000001n V_low
+ 998.100000n V_low
+ 998.100001n V_low
+ 998.200000n V_low
+ 998.200001n V_low
+ 998.300000n V_low
+ 998.300001n V_low
+ 998.400000n V_low
+ 998.400001n V_low
+ 998.500000n V_low
+ 998.500001n V_low
+ 998.600000n V_low
+ 998.600001n V_low
+ 998.700000n V_low
+ 998.700001n V_low
+ 998.800000n V_low
+ 998.800001n V_low
+ 998.900000n V_low
+ 998.900001n V_low
+ 999.000000n V_low
+ 999.000001n V_hig
+ 999.100000n V_hig
+ 999.100001n V_hig
+ 999.200000n V_hig
+ 999.200001n V_hig
+ 999.300000n V_hig
+ 999.300001n V_hig
+ 999.400000n V_hig
+ 999.400001n V_hig
+ 999.500000n V_hig
+ 999.500001n V_hig
+ 999.600000n V_hig
+ 999.600001n V_hig
+ 999.700000n V_hig
+ 999.700001n V_hig
+ 999.800000n V_hig
+ 999.800001n V_hig
+ 999.900000n V_hig
+ 999.900001n V_hig
+ 1000.000000n V_hig
+ 
.END
